// MODULE : VFPCONFIGDUT
module vfpConfigd5mCameraDut(d5m_camera_if.ConfigMaster d5m_camera_vif);
import generic_pack::*;  
    VFP_v1_0                  #(
    .revision_number           ( revision_number            ),
    .C_rgb_m_axis_TDATA_WIDTH  ( C_rgb_m_axis_TDATA_WIDTH   ),
    .C_rgb_m_axis_START_COUNT  ( C_rgb_m_axis_START_COUNT   ),
    .C_rgb_s_axis_TDATA_WIDTH  ( C_rgb_s_axis_TDATA_WIDTH   ),
    .C_m_axis_mm2s_TDATA_WIDTH ( C_m_axis_mm2s_TDATA_WIDTH  ),
    .C_m_axis_mm2s_START_COUNT ( C_m_axis_mm2s_START_COUNT  ),
    .C_vfpConfig_DATA_WIDTH    ( C_vfpConfig_DATA_WIDTH     ),
    .C_vfpConfig_ADDR_WIDTH    ( C_vfpConfig_ADDR_WIDTH     ),
    .conf_data_width           ( conf_data_width            ),
    .conf_addr_width           ( conf_addr_width            ),
    .i_data_width              ( i_data_width               ),
    .s_data_width              ( s_data_width               ),
    .b_data_width              ( b_data_width               ),
    .i_precision               ( i_precision                ),
    .i_full_range              ( i_full_range               ),
    .img_width                 ( img_width                  ),
    .dataWidth                 ( dataWidth                  ))
    dutVFP_v1Inst              (
    //d5m input
    .pixclk                    (d5m_camera_vif.pixclk        ),//(d5m_camera_vif.ACLK   ),
    .ifval                     (d5m_camera_vif.ifval         ),//(d5m_camera_vif.ARESETN),
    .ilval                     (d5m_camera_vif.ilval         ),//(d5m_camera_vif.AWADDR ),
    .idata                     (d5m_camera_vif.idata         ),//(d5m_camera_vif.AWPROT ),
    //tx channel
    .rgb_m_axis_aclk           (d5m_camera_vif.pixclk        ),
    .rgb_m_axis_aresetn        (d5m_camera_vif.reset         ),
    .rgb_m_axis_tready         (                             ),//(axi4l_vif.AWADDR ),
    .rgb_m_axis_tvalid         (                             ),//(axi4l_vif.AWPROT ),
    .rgb_m_axis_tlast          (                             ),//(axi4l_vif.AWVALID),
    .rgb_m_axis_tuser          (                             ),//(axi4l_vif.AWREADY),
    .rgb_m_axis_tdata          (                             ),//(axi4l_vif.WDATA  ),
    //rx channel               
    .rgb_s_axis_aclk           (d5m_camera_vif.pixclk        ),
    .rgb_s_axis_aresetn        (d5m_camera_vif.reset         ),
    .rgb_s_axis_tready         (                             ),
    .rgb_s_axis_tvalid         (                             ),
    .rgb_s_axis_tlast          (                             ),
    .rgb_s_axis_tuser          (                             ),
    .rgb_s_axis_tdata          (                             ),
    //destination channel                                    
    .m_axis_mm2s_aclk          (d5m_camera_vif.pixclk        ),
    .m_axis_mm2s_aresetn       (d5m_camera_vif.reset         ),
    .m_axis_mm2s_tready        (                             ),//(axi4l_vif.AWADDR ),
    .m_axis_mm2s_tvalid        (                             ),//(axi4l_vif.AWPROT ),
    .m_axis_mm2s_tuser         (                             ),//(axi4l_vif.AWVALID),
    .m_axis_mm2s_tlast         (                             ),//(axi4l_vif.AWREADY),
    .m_axis_mm2s_tdata         (                             ),//(axi4l_vif.WDATA  ),
    .m_axis_mm2s_tkeep         (                             ),//(axi4l_vif.AWPROT ),
    .m_axis_mm2s_tstrb         (                             ),//(axi4l_vif.AWVALID),
    .m_axis_mm2s_tid           (                             ),//(axi4l_vif.AWREADY),
    .m_axis_mm2s_tdest         (                             ),//(axi4l_vif.WDATA  ),
    //video configuration      
    .vfpconfig_aclk            (d5m_camera_vif.pixclk        ),
    .vfpconfig_aresetn         (d5m_camera_vif.reset         ),
    .vfpconfig_awaddr          (                             ),
    .vfpconfig_awprot          (                             ),
    .vfpconfig_awvalid         (                             ),
    .vfpconfig_awready         (                             ),
    .vfpconfig_wdata           (                             ),
    .vfpconfig_wstrb           (                             ),
    .vfpconfig_wvalid          (                             ),
    .vfpconfig_wready          (                             ),
    .vfpconfig_bresp           (                             ),
    .vfpconfig_bvalid          (                             ),
    .vfpconfig_bready          (                             ),
    .vfpconfig_araddr          (                             ),
    .vfpconfig_arprot          (                             ),
    .vfpconfig_arvalid         (                             ),
    .vfpconfig_arready         (                             ),
    .vfpconfig_rdata           (                             ),
    .vfpconfig_rresp           (                             ),
    .vfpconfig_rvalid          (                             ),
    .vfpconfig_rready          (                             ));
endmodule: vfpConfigd5mCameraDut