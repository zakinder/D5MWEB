// MODULE : VFPCONFIGDUT
module vfpConfigAxi4sDut(axi4s_if.rx_channel axi4s_vif);
import generic_pack::*;  
    VFP_v1_0                  #(
    .revision_number           ( revision_number            ),
    .C_rgb_m_axis_TDATA_WIDTH  ( C_rgb_m_axis_TDATA_WIDTH   ),
    .C_rgb_m_axis_START_COUNT  ( C_rgb_m_axis_START_COUNT   ),
    .C_rgb_s_axis_TDATA_WIDTH  ( C_rgb_s_axis_TDATA_WIDTH   ),
    .C_m_axis_mm2s_TDATA_WIDTH ( C_m_axis_mm2s_TDATA_WIDTH  ),
    .C_m_axis_mm2s_START_COUNT ( C_m_axis_mm2s_START_COUNT  ),
    .C_vfpConfig_DATA_WIDTH    ( C_vfpConfig_DATA_WIDTH     ),
    .C_vfpConfig_ADDR_WIDTH    ( C_vfpConfig_ADDR_WIDTH     ),
    .conf_data_width           ( conf_data_width            ),
    .conf_addr_width           ( conf_addr_width            ),
    .i_data_width              ( i_data_width               ),
    .s_data_width              ( s_data_width               ),
    .b_data_width              ( b_data_width               ),
    .i_precision               ( i_precision                ),
    .i_full_range              ( i_full_range               ),
    .img_width                 ( img_width                  ),
    .dataWidth                 ( dataWidth                  ))
    dutVFP_v1Inst              (
    //d5m input
    .pixclk                    (                             ),//(axi4l_vif.ACLK   ),
    .ifval                     (                             ),//(axi4l_vif.ARESETN),
    .ilval                     (                             ),//(axi4l_vif.AWADDR ),
    .idata                     (                             ),//(axi4l_vif.AWPROT ),
    //tx channel
    .rgb_m_axis_aclk           (axi4s_vif.ACLK               ),
    .rgb_m_axis_aresetn        (axi4s_vif.ARESET_N           ),
    .rgb_m_axis_tready         (                             ),//(axi4l_vif.AWADDR ),
    .rgb_m_axis_tvalid         (                             ),//(axi4l_vif.AWPROT ),
    .rgb_m_axis_tlast          (                             ),//(axi4l_vif.AWVALID),
    .rgb_m_axis_tuser          (                             ),//(axi4l_vif.AWREADY),
    .rgb_m_axis_tdata          (                             ),//(axi4l_vif.WDATA  ),
    //rx channel               
    .rgb_s_axis_aclk           (axi4s_vif.ACLK               ),
    .rgb_s_axis_aresetn        (axi4s_vif.ARESET_N           ),
    .rgb_s_axis_tready         (axi4s_vif.TREADY             ),
    .rgb_s_axis_tvalid         (axi4s_vif.TVALID             ),
    .rgb_s_axis_tlast          (axi4s_vif.TLAST              ),
    .rgb_s_axis_tuser          (axi4s_vif.TUSER              ),
    .rgb_s_axis_tdata          (axi4s_vif.TDATA              ),
    //destination channel                                    
    .m_axis_mm2s_aclk          (axi4s_vif.ACLK               ),
    .m_axis_mm2s_aresetn       (axi4s_vif.ARESET_N           ),
    .m_axis_mm2s_tready        (                             ),//(axi4l_vif.AWADDR ),
    .m_axis_mm2s_tvalid        (                             ),//(axi4l_vif.AWPROT ),
    .m_axis_mm2s_tuser         (                             ),//(axi4l_vif.AWVALID),
    .m_axis_mm2s_tlast         (                             ),//(axi4l_vif.AWREADY),
    .m_axis_mm2s_tdata         (                             ),//(axi4l_vif.WDATA  ),
    .m_axis_mm2s_tkeep         (                             ),//(axi4l_vif.AWPROT ),
    .m_axis_mm2s_tstrb         (                             ),//(axi4l_vif.AWVALID),
    .m_axis_mm2s_tid           (                             ),//(axi4l_vif.AWREADY),
    .m_axis_mm2s_tdest         (                             ),//(axi4l_vif.WDATA  ),
    //video configuration      
    .vfpconfig_aclk            (axi4s_vif.ACLK               ),
    .vfpconfig_aresetn         (axi4s_vif.ARESET_N           ),
    .vfpconfig_awaddr          (                             ),
    .vfpconfig_awprot          (                             ),
    .vfpconfig_awvalid         (                             ),
    .vfpconfig_awready         (                             ),
    .vfpconfig_wdata           (                             ),
    .vfpconfig_wstrb           (                             ),
    .vfpconfig_wvalid          (                             ),
    .vfpconfig_wready          (                             ),
    .vfpconfig_bresp           (                             ),
    .vfpconfig_bvalid          (                             ),
    .vfpconfig_bready          (                             ),
    .vfpconfig_araddr          (                             ),
    .vfpconfig_arprot          (                             ),
    .vfpconfig_arvalid         (                             ),
    .vfpconfig_arready         (                             ),
    .vfpconfig_rdata           (                             ),
    .vfpconfig_rresp           (                             ),
    .vfpconfig_rvalid          (                             ),
    .vfpconfig_rready          (                             ));
endmodule: vfpConfigAxi4sDut