  `include "../../agent/rgb_agent_pkg.sv"
package rgb_pkg;
  import rgb_agent_pkg::*;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "../../defin_lib.svh"
  `include "rgb_env.sv"
  `include "../../test/rgb/rgb_test.sv"
endpackage:rgb_pkg