package axi_lite_agent_pkg;
  `include "../defin_lib.svh"
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "transaction/axi_lite_transaction.svh"
  `include "sequence/axi_lite_sequence.svh"
  `include "configuration/axi_lite_config.svh"
  `include "driver/axi_lite_driver.svh"
  `include "monitor/axi_lite_monitor.svh"
  `include "coverage/axi_lite_coverage.svh"
  `include "axi_lite_agent.svh"
endpackage:axi_lite_agent_pkg