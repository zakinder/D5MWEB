  `include "../../agent/axi_lite_agent_pkg.sv"
package axi4_lite_pkg;
  import axi_lite_agent_pkg::*;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "../../defin_lib.svh"
  `include "axi4_lite_env.sv"
  `include "../../test/axi4_lite/axi_lite_test.sv"
endpackage:axi4_lite_pkg
