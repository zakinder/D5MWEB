`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
WSNqUWyxzStdcAcjzmbg144gkTI5BCUVrPWAD5aOuDNiLLteNB6KhcQLoE7OcCCj8Guuu1xncYvu
Bk8rkEJtMQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EMRgPNCcrZHHKbd8g35GpCj96pJM85AYIvQE1eogue2SjS7tKcH3f2cqc6dskKbmBws+qZjVZM6c
h7j9CX8H3V73Yjlblp9QuD3k41FvfBdz3Hyc1Vgh6vaLoW7MCt1GOREU09fH8IIYZ4UBGMWgDjXM
xV/TNvV5Gv8xw+h8cVY=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uZKEDXKcEzzdPwDayteGLiYNYbrUjcl1kd3JWyM/Lhm+OLhF3b2mAr9DcM4Zazc48xCTHRT3YMLu
QugNL8D/i5mg5XgXlIR3+qdv11PXVV6dS+XNC4uUoUcJGxIrVTY/ZS+p/kGBYrZIo1YdSDjcMubD
44CcQp+w/btfIgQGQIY=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
x1f3fuXklazmiiEmkGHsbEIMKKFZZKbSvAjsHf+Fg9ED1WDA5EM29ScXH4/d23JW0hyJf/qKGMEI
amH+QeMJuuaNXaRispQ/5BUoWup+uPqE8X3lvWPQUaBoImwv1rdVChAK5b19ElEDFpaKXnpwNA+t
ORC7Z6cRKe7He/k/UM2PkeoV8nq6HJX1dU/6sQD5PuAC85dAOhwaaW7GZ4T+nsFCTVmcE7tXXIaC
v7/odO3RoPmwika3IgHSqdE+8hyAgXShOAFT/16YxymdYWU/j9Gh/DB23i9Gy8ZzDmNczfygywPy
wd3ojeyMT/qaJMDabt1UJ116r4GhNAnqDSRmbA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Zol7oY7c/Ggo6jliVSbanJud3kxI3TGEJStU6oh+w207/84Utk4j3fLReVcx6hDQ9Y36Bde93klR
zxdGuusXOCmcV+xazZVNxqYOvoC8nsG9ZVomATSFgyWYJ7MzQBi6WsjR9tG93jH33/RmMhEjw1Od
J59qm2BBpQz1dVmBFYgYBgGN4NKXeYkVsZTBeqCYh8OhFPitnrszPEJ/JLREO7JclKbDI8BY46z+
ON2Uly6M39msk8Sz7eqSIf7UGiMcHhcuyFbex2LHwjN9OJjHY9NeWd40ZT1NXkCJWgEKHN3T4tWJ
dTpGvezqCsdVZQRy6/KLkwXaXjsuiPzfMqggKg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rlO7EOXjAX98xk5WgJRV3KPFqxeNdX6ooTM5jCcC3CxznQ2ZyjUO43H8J9pXrkzDLjBX3eVTI0s+
Sibzu7B8XvJAM+Nl01WsysdGLAm0npS9Cn3+97DjCt5QRxJJFzNlZ7FCYQn6pWrDypl2Mv8pmPWV
oBFRYsjLGOZ1O/1puMY3rHiMb8bPSpkS0TDh+wI4vWopTFm8Kj1+LZCHmvqMFUVM2MtmElCBq5bu
uLFott8WIilsd7UEXBh2DhQiPQSN0LkVj9yk8rkz4FAigGihoxMhyQAxufO4+t9dSq7buFUUEWwa
OYeETiPq9EU3eQ8L8Y95WrHebWXeTh5fdD8LhQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 63104)
`protect data_block
bC2+fyeM27+JMZWyelQ1uUpBeyqlmgLFoyS2RxGWarSJaZWyn+yBXbZuMokVaHLuo0qxPyMWr4qV
uArDQYwpVI2EKMl7PurGPJEjUh5q3F6oLgOBWWyHcqLmU0XUTzfOBLCrcRy6+CkGYrezt0s9M6kr
k4yELk+jUtye1IVkdm4q+rlE1CAwPQR0T7eHHoyvdAFB1jfX0lF/DvsRulGMWgk5h66i08sgZFif
Kx5UqjvASvgGaZDZpDZpAqH8iG8KyXjGnvB84YkgD92nZGRIh/hsxMfquvZztBEq4OeE8X9DqJSE
w2sswlOJm38AjQ8nSfL+b2m3nBYlii0E+5q6gXkdv+jIrTwuIsLYs+QxYKJLaUsFiefe8SYYBXrH
JjZPqfWTMy9UC+S0QBeqK+BjoJVFwl61s5XhBGUVe5k9SNgvH2j2E0f8B/4qS7k8FqB1FH2uw7Mx
BvQreTzDlhylAMwkIWYbZqaHwNP/DwAzSCwjfvIgDwpptUdBo+EArarqgJKMdQmZZ3iNsDGH3GCF
tyeZglwGr20v2HNoTVaJu9YsWm3qaJ59VdDJAZ9FGAp7hjiSOBvtdNNeYA/PFQRUVQ4w3UTXMQ0d
tSaWLUfhxsOe4poy3XB9e7VSCBOXXRjvNfqa0zn5iOyIUHWNOIUrOlejeMO/UabF58aIGGn83qBU
NTrIEtw54hqB9p0kl/syXy/DwigE6b1xRcdYzx8h5YmyV+ZRDqb6biAU3OWybHUQuzlEMQe9GW9+
D6sxeky2SeeDGkHnUgF1sgnrQmZxOKAj6fK1pIiIjHdpdv+FQPdG5ienaii1y8glBvfVcqg7G9kr
rnDlVduPoYLZOos0uevDR5pa4YKk2eEXzYd0ObbtFVxTA6dC6yMd71fVbhNRP5DR27ex1XlaNCrO
gOD2crOAVYENJcXFKMKoKyUfjzxvyq06gmfPMRVJEqWjNmuRkArjfqY74NCEqMwHIcjFU1eGymvM
2UcWs8P0haPy6gmDl9QKOhXH/2dDM4gelzqUvg8yB8m3VDKZY8fPN898bmomZSaA/l3eUIMGt8cS
r3QBEJ7RwRnlDBNS5gAAEKxl9TqK3ZdaK4O/c01LNjj9p0XMH3LX7E6Jt9CGoizoWHrMO/buYF7R
Hx4ubmIWWj3rlZTD77uM2RNJUPlRtk35Os+Qp3wrHDSs5yNQDTbw0OYZA9V0w8nilCfGQrEyZOQG
xzYzd3yvRQ2GfLVSkjE8bjwZCS3oQr56uBfuyiuBfeK8utD4LdTu4RevNaYzfdX/Ct/A/nHzMRtH
4J0gJ0YI5GjMT+BShiGxeShC/orcdFE18geb4fEODXSSNpTQbUqhJNXW3i3frdZxZp3tTSiguaw4
jArP5jlbzQmIaGnb5622Lyy5l6Lg5jW/o2is0KC0LvTACMfyRO4cpSbEPRpXnXsA3GbS03Hgsesw
/HcelQvR5gWpJug6/VXVpKPQtkkVTKIND4KhLMz2vixfUNwT6VtyHnhqIZ1zcjVh0tYJ6BAEaC6z
vUCtz41l0YPVdvbMrJDr9GMbb/6PFn7h3qm3gzl10+xzJ5mgEwe8hZ6G25ksSK7r0Aewlovu6aDg
Vv4Gcd8EVbGXsnOg08lqBxBgh3e3rtMFvil4pITtpj/yqPg4fY/unptTwDeKZ91aLqhgFXnMaNre
c8uK0qGqFsYBl0pwywKH+kZPP3m+K0QqOgmeMV1J/nOzAmOKDYa7ksZFcQ5fJMPWjk0q5SqzV+z1
Jx3PRYAV8OlRQCWUhstdNPrYL/Y7x3XbE9+Kk9pgr73lRnoc8tSNmWWpip4l5jR7IJAkZ3iPX3h4
FdD9J/zJaBniQmA9RHCb5iOuZdXTg2CB2+mCk9qYZ9yYllbvjVjip1xltCMg1rRfdiO2d6gnc4cM
rmoH+/LCCwR0XHkWP2P/IM8dlFuF9ZGqk/KavfyPb8RAPOTkrMRynP4ettxXTDsHkvJtdX3B8BdQ
d7RWu2kLFkLMfM8DDSg26KgmvjlNBfvjAfDLgel6Lmm/ZI0KvPLoX2t4YMNNdTVVTT4h3FkaJPFZ
+roENqwx3ChBuF2LsjouvO9nCiHy/THdqMxKtWhawjmQDEjoh2XUAXQKa9ShGBK71oHTNTnARwDS
g4D1LC2LcLAsGSbwBl3X4Nw5pZKiPJFPAmYPMmBXMIwclj6O0oB7ktF4ae/pwCmasirwQFO1Yceo
8sJgdhr8AID8+eWfu+7nblMFGgk0PzUskmRJp4rT+v9U4PbqnYfPQLcZnofTqnQkT/9wTcAf7JMk
3ZMt4ns6Ku6yzzM/4OQqQluo5Te7Onv2CuYhiFYFFWaahdz3RfNnkJEF1kCqwtxoG287tC3ydH4p
9LQdKa/P8I5Xcmo5QgzUep353OGsaUcwgisKrBwv8PPAaIpVC+d8xn3aY28pGwLerchANprrPV6y
yctu2BBdQUKK2zRYr6dNM+hoI+JRrsWUuHPru5yxZYMUEYzf5Kdw1evFzU2P2PCdn0p4ScVORSgP
AblOf7sb3xvvA4aJssj6RMvM+WLjxqtP3qenI6AKh+fZsRGNxKYjKcLJoBnakCXr6N0EWuwqWKLO
QPyue9AS4JhHuFlI+hxRkftCzoTKS8ZgI8LKPewdvw1kUHINlb18zs02BdIQ6jTLQi+bD1y1uo0P
w22TVabBqEfxpFoN3GvpzEb/bWoIe1GcakyfKa3N857afnYkAMTULEK8K9Q09h/Qt/3zX0S0uVO/
NDeFWzEiJoC4Uo/jOY1at/4Oz2oREERP8HTVRh1QFvPxyULVUO5sWvMbkhb8HS4N5DZCsqHtoHf/
G7VEC7ojHQq5YJEPGX5LuAD9KOy/fHvyYhlp7BwXgaBfwWrJ9/3BM4z3i+gRjxxL0OhenRZiqtpb
uINYQUjVX3LbePo0fmcXQGVrDbIRANauRIedD36dZ4n7WLn4IDKtLC12IOABSuDo/8KyxYBKFDES
rB/A2c0a4l8D9nUyvyproA5hkctgn9csINMdlVrNG3R8/t+QB+2JFP+AjcuFkKJ+KedNldC+Vbiv
d9VnEfubdkSXgBun42YdTLGL9/9w/H+YUkByk1W6VJKk9fZ0daYWoFdkMKL98Pje5zi01sCdLNuE
n0wUGwQX2l5ChCFwRPefz0Ckx/S2TjnhWqD1eAb6WVh67vchBraEO5fm5f1bp2zO4NDTsND752Pk
OOj3oVJSBLJdlZcHhxDwMxMGJOd6U0qudNdQZ+i28wMyC7yzyDJe/oYbgLYMav5dGu3hbTOmGe0s
IOnw/2TRpbxpt5ofLw797yBvMBIdMBPjnrln9bfkBCDbLHRJxamoLa6q64ppPyL0MZciwrW9r+RH
EOKFZshB7l1poKJvTon2JdAMF0+1ul1pMhNRcCaj/F8IWHpilMOEntkKomnhBmtxypriSObSOjBo
/B7rr/IegyNwCaSipIpPi5P1cvrTTVTDs+tuXWqlunXbMZBsCKmVhQ5XLosTr/fYYjyitVIMlxGW
1KxFo2faUNoVufBXHzD//2d3zXde2guR2r4QpDU38cHpusTjVL0isj7M4ZSwuzDf2VR80eFIgsrM
AW1oV+MDUy3wdBYDb7ZDT2TMOAPmatZ92EF45Sol/EneUuLyPrKr6U8wV1kzlecYHr9PB3uQ5NUF
7M67TiPb45+j9TJXTJo/YO3UsTyEodasWcAcabghuJHRNew/4nywqUhjfr/e3w6JCR3oMDXLYzDx
WyHfw9H14RxwlEMiScVlF4OYSWsksjp1tUhgLnn2NXPks2pXjLacQ3uKbjxXcREaJiOIJhV/rBd1
M1ltQZyB1mU/OTTf28a1lTVz9VR7QC5u7PKtdS1XHaSI4EiNNjYfzBz/QhMCcJMY4Peh1N4SavPh
J6ZSQeXLmVgedcLCN4Yj5x4nPH7lQpcqlXD833nXZPsx7ZzXIOBrjSsS0yNk5xvL7gsldjdRHTHP
6QL2iN81z/5SqDAlQHsJi4Zyj+FOuvJyViVdQS1RXSJr8M5POPeqeYHiJk0JjwYsQKMGy5IRtdy4
lYNqlmwNPDcdBt+AkI+xPdC39E6AqrEdQGnYrNJ0NRW8yMH9ppqadA3OlldXRnutHxVxq7yqKeWQ
XK1SHTZUi2MYyJOetFrwiM3h9AwPeiLK6/k61A489RrGZiBVqo0YT9mM1qA2QrkXLD9iEGy5ydcU
sk4jHNFc2wO7voezrU2M+RDEFxxJGDSoIVwaTvyHh0XMJq/Qs+E5zzylK082oLDLJvxBub81Z1RL
sKRK3tY+70jHfRtOaecGSpejRVSrmvVZrLEnkJtPud349gYlPmeYEKwcNlncVRyr0yBqrxoCQ+Hp
W7s4lt8ZUdAGd88fbEb3nYeYUPSsZLx1l67VcXjlsO6knopNftdzLBZArvZWUk88vEaYOzpfy4Rr
EQ14qjQ44r3Q2238CzaCtzuHX62hj8o1N0PhggyQZw35LiED7T9WcxVZaVIhvBRDRqayVu7bYt6B
gqophIwmIdOgY2tN3/B1Nou6ApQdW2TaCnXJgC5JHySW8yfphfohU1+tLp0gMrNMd5iHGbE446C2
BDEfHpqBjQXn38P1mYDJ8GF3N9Elb2ZHGZ+rbkv2qgy3oAcIh2DSkyQ+DoFx0NXUMmx+so7w/o3+
IqdX8MT9rsT55uS509EhhS2LMLL+p3B332+YFqpmorjW4djfmi86R6r9xp9FuHj3c2/oYLUu1aLq
zdW5lbLShHZ4M/FB4nlNJqbThTLGd5BJCsvnzvN9qeENkCSB7DJTfdT5NI0OW173kMdmmmqv4VIs
gui6zbUdQr2ffJ91rkXq7aC6y1/Vrce4FXOfCRt4oiwkUgpqQvHffX/nPMsPC1mEb3MlUbhsjqeQ
Utw+UgR8+7ulHSX5fPfpBTFtAdxg0iLOdBFywE5Y805h9BZZ7/f8BU4sOQyP0GECDwhkl9b/doA2
JwjgjV1XRyhzDVmwZVvX1c8EMwyMdTuti3HszPKaVNMYre6RnfDsJDWAaZzIC/xwvk+Qc5i6XAtG
5knYLC6FYOtKvMFn66gLq8xMed6CfliN0fYLAf7I/+Jh8N+jb+Lit4a2iH/iwL28MF9FEXbPGGNQ
vvztidBigyLYuz55juNSKNPv4LfId1gM3p/Ph0hVAWnMdmjsFJgB+ZfHy7zYtdjcRw6Nw0LXzmku
XVcgVr6ozDGA3fAzJPLoUeRqr+bStE+wS5DEUICPR/eO95zIoMVzgkizJ1fiUOaAkgRmXkdQuia7
yEpji51GPfJROd5Xsa0mK5VFnrV+N8XWDEbY4Xks32HfN2ducoTLsS4lIRFHaTgsjFHdO3RasPUu
qjAqFbNO9tgonD7gFYbtYSv9qLBEufDmSqOBPgjJRMGWTzyuJI5vaQGUe5SdhKI2VXxK1cgLZrI9
+C/pTPCVJiIcEHLfjMKCla3BzbMuKMbTv+Uag/lqLmf5hNDesw2qoWOh8kr8fEBvDDQVHHt2xSSs
0IN134lEwmKQlMnYAaCAK7br3s5nm04YpfyaBYSa8tP50nD4MR6Wa73TkP2CisRW2AO6XnyA+xoN
TO2vjHspYR8HBLCRjcjvebaG9c2/Q7ouKqqPrhSEM24CfQhB1gRc5Yp3WjluLNyWbmWU8KNtRoP2
8hF4ZFDsUnwZ2msIHGuLO5O9ZZD7VFPC0JyNmq/D4zB7REY5cmt+WcP/uNj+zJ133PNX8JLwkHnk
oKSkhNwXfTe2IJjuz6evl3oNtsP/qh/NkEZ11ONOebHP/JpERkIYA73gLP+NMfZuYHmUHf8PXXO9
0deCyK5ztLfQ1j1UTZM5rftB/sRPy5DXK5ROMUGCjS61xkb+S4iTbJyRA9lTawnzF4/pLvdYuYhg
BVgAd8RAodn5EVq4JNLtQxPKKni4qKR8nOGHZGpJVkk/e8qY8J2r2zh/Xk/hSMZ8uVZyS+Y122Ru
+NXBNczKNH7Pwiwjls9eiljx2OrUKKrE9cIbtUSLrnOhOdi4QXbsw3xix0YaPJMLXLSPiVYIC6IJ
LLH81hZ1KS2b8vjHFItu9mKZbrAB5FVBssoHpKcnWw6bv9+IEEORY5E2PaV8t0vEQALchMep2hxc
xGs6H9/tngfHKKEmGZQyFG9so8rRziqcMu3Edr8Fj/hTK8Tcelvrz9NpGKP3/t6JUUctkk/hGa1H
Ck5c9Rz/RzA23vsdhMkHTP4GMyrRfk5LUxoHqDyOKM+W5czbL7Hzw5/Zt/utRvXYP3KnoI6h0Gm4
5CcRo8ex4P2e3ET4dZ0fHsvaM9TBtP+bzzDXbc0TLaw90G5Gz2nEORLyYzKQwREzuN1Y3cLvs3Fm
1clEt9igPsiFVg35hbOeTBQlw9UftCxxec4H+jNv20AiLCiXmBGAzPu5T0ETZ1pN9Vgj7A6hcBrg
ENz/Fwqf9npnAe2wonXeZYxmc0qKElwiybbWY8ONcI1XUmVrVVPzuq/DDLPMnWF/NSfC4dDst8Ls
6iv1Fmi69JV5MhhEWf5wIvCYrs4k8S052u4xHGl1UzDCG19O0hkIU7VaneVeHwOP0kOyjy+AqJY4
z0DuHFNWi0+k+Smd40u9Fke4Vkd+vsadkt7p+tYVMN8xzI0gNlgoWB8K0xIuEg8iqITNtvOvq0CU
I0DoKkZsCfOwCE40hZgeTitr5dQCe3xk4CDdJQWa6mePutSKM+J8tGpR1xUf5pkEw7SiL7H+bWwT
uivAdxYZqSZiXau4/iutRt6V/NacmgISUTnyM6LEY1Bb8T6y17UFg70H2+DrvIn3rSTmJ68+fN9i
YwyxHmTV7RATxFSbovBrTVRSESHroPUO7j5Q3kZtnADrcWgGXHHbH2wsKVPuMfZFVIuh1eIyZ01q
sDr/qekNPvhC1j4Q0vHQdJ/tytZMeaxPRDmWyUy1YclkIKVVR/jVoO7KcoHNxXebvbgFwgtNdud7
qnWdYAOOEBul8IGqHTXJ4Z59LJtmwK3r6xDRGxSnKfpK2zrt21w1bblKIT/QZ6TwFkBNHjZHyLnL
Mycmxt9pwSwdoscM/UdqqDGE5Er+5CbIWSywmdcAum23O2eoWveow05mepDoeVl/zPYuPdNUV9+u
P/TRknYVXXNuDs59AvMKbD/Wfe6TDI8nO67zwR9UQx9P0Ra6hJyvkZUIo6HtVedJ9XQ4WqYVIUzE
QzvAakLsCb1XQPvFsBN5006q2/An+eTY9QVfcGc6NR/pEFyRUHK9fgC4e9A0uLnkh/S/TDYK6Jc4
CrPRhFgm1UI7thHH86XXLi+JZ9n8MZiMhx9NmrYVsISOVPD6dn/cBsLOkMYEfPCHZjx/Pn8OL+42
KmPyiaYeLr3MVPUriMFbrvMuBeyzvAn2jr8THpkQ4GaXR9nUTDrN7Of4bC4cTu5xbHJc2y4uzwTG
WT3QWDiuL4Ikc05DUXxGyniMPgmzLC5Mf4D1nqImSktvhIoaUHHgNBY/LDXK3ZIvjBrDNcqZANNR
lIWvGH7CN8OOQ3Z6uOzYtm0yWuetqfRWiL9X/sSqKEgwmi3miUVs3I5H7Cm2HpsO/qBc4Deqda7g
D15NEtxCA/xMgM2clHXTWflXwlkx0e24afhXBl1LtmzkfEwLbRBSALaCgagi+IUY8mnahc+GOCC8
Yns8DUFcsDORl28Obk8n7ZW3wW6GcQMNf+2J95L/crZlrk5OL1BXCAkfaPybgPRp28cB9tP/I2TZ
y9aUn8ydM5d0j9qCid3+C+Uuhmc1eaI7BQILyM9QHoD/5J6CmhiIhs7WMefXlGjhjN6DpPJNcmcd
a65NmejKZIJDQY3gDu8w7pEFxolpWOulJXAF8sa1uGa2PJAaGCoV60nkEYAN3tHBkh12at7TgMAA
Ad0bPfY/5zM80KPzKFKDNDkQvsp8eldxuf5ofLsF3LI40Tiq+q2ATVV/iOq2u2EcynhuTbXziYkn
tiOKypNC9dOXugME5wIKQ2rEu6va8eC+lP5hMa4ETgU0UNVSFp7v9AA3170UiEYyr33dTItqnBR2
IEfIv4g6prqK6OQHJh863EUcJLkhf5HYn3u3bTBC2fSjQyQ/wn8he1uiyp08eD4w7zNg/zuH1Jfu
9dsEKsyv+baiS9iTbgzZU8pLenbqUqxx2Imux+/eWvTnkod+gjLBJJ3OaOgCSj53ARoylpvWmnYK
JD0zCWjYkS/qciLRq1KLeUyPnI1XfjfkJO/8vVRKjHSYwnIYHtvZ/UrfwLnRXxsFSBQQ/vJXy9nd
n9LPSwvSmV4eSxQhv+2DIwlsRxdlTPm6sUTRQ6C04mg/VkNXtmqGEcMJFCHbS0mg5/g0OKSe8ynS
1LrqLWilEMKTlwb6S4aWcPJ7MqVoMLqE4ICfoI71XJOIYrxK2UQx1LmNcsFgEVFAU1cqqWXFJw1w
3atO/rkmtT3gePAU/HYA3YYBLdWGpEt1qi03rs1izoxGNC5IRsC1drfms5zBJLfQ9mBZhUHVtwwQ
t4hQh8FRDWCV7LdjA+temtUeTWmewOV0/OXAK9RVsFFD3tbi1b4aW4jDhd5eDOIQgYIeexLroPkU
nrYQgbgtJP3d28CGa/upbnBGiQ8hAF2SfRmPHeQkXssR4fdCGXk2+hp3icX789XXKbGlic0ex2uI
EcZuyDGsvJiddCMII4gW2CuSlebhh3QoH6Uol2KA99WbxGkXecfo5BLv15MATtSfqZzXTP5RyR9w
AwosNyTjaokrQcKnTZlzLP84TjGcGp2yKShIy/00OgMbgLeCuKPHyPCZSsYvgd0alxlTVrWRXmyi
ASkZz/7kGH9sWQfGV4I09OMIVFYn+Ub9GO4D9Wi+XOI5ipTYvLn1s3QNNZqcf6HKm/eUaUDsKkCY
3WK5kx/8qNNYkkeYVs3UewQov4K5lw1AVqrXd65ITPjKEKj3TY6VRE7GwLyvdJz8RBN89FqKSk46
iNebxKQQ8L6iBhY5c2L8yQvKBCe2pjprtkEthURufD2Y5NaRjYBVS0i2ufjpeFju+bu6JC1gp6zE
RmjYJzVoZ1OoHNckGZ8kLW8aEQZvM+Qw0TUEFmPQfjvHgRcNmUiGFpMZlAmLFHZE2w/+SQqqP+kU
55056sx0LO8j0POssjLto7OU7bL0/3DbQQzeYWpKRkKzsvPn8/aMUmycYjqAYUyGxUzeCn2dUdpu
b3VZhME8Pg3Y963tzR4YhICNwjPNjdVL8J6fy9703SGbZDWjWw9LbkQwlMYbKv6vaP8Aipcoqk5K
AljoJtWA6a95WiqQZPKH+rnrwJ2Mu5d/vv4Yz5IWjoVzEIyQoTcTsu7nNy8Ip998AttMb9P5323z
78xslK6iNIF0X+fq+fvkqtrQFDm568FPJMkEX+ekAP0WHK5mi1t1GGHPzB2oUVFVgQN7VauySq0g
Z6uCc+AqJNBnAMoIehtcPe96ox4Rwq2o01rgeb3DDGq2S4GdTzLavULFWMc00UPVuwnuplDHEyNs
/AcU872vO0Leei+tl1pSwQs1wwDsKAO+FUQkfcW0SrCm4YKmB7XlDfcQeFwosIA9dXodEHkczGDy
Mo1DMRJaAPa0L0X9e0aGkrjLoX/9upVzhON8wBRsGrzEDLVpTIvy2aPDGVNV5tOetMr7J+jhimEO
XRTgEeqNv8kbyazLL5WJQI3B1EWqUqiP5/hLKp4sjHnNQ7yjDZnw5CoomdnEfRByOTuMxnHc9KvT
J8N1+nEBDnd1TM2fdu0+cSFNW0/1j24Cqr6pfacA4/AfdNUjXU2w6LHiZE5zIKD+Yb6Lp0jkIxzj
JMJUFmO6VrgQ+W7n7lYc9H2sctbe1lWERRDWYJY6cbiXo/x7R2ei/+uu4QkJscgXLO3ifGBA9a1B
/rn8Ghpq//ZRekVUQ2b0x2GljPIqN7fY04cM/gfPpzYOOFvQS1IqJ0r9sulI9vbwxGBwCi4l7Jbh
xmDFhO24vosOIo3n6yUyxDbrqsC1iqP3GzKJ+Aez4jsmtgNOsHhZo05N3rOAwQknKW0USs4xVKpp
px2Fdpv2xwG3tNuJHJJOLdDnI5JLonFSnCArz8mG1uPLi21VO55G07HwgxC4tEXbu85CRDmb5pOA
OybGxLsg+LLNFGyepu+Bx/bpYQ4gam9ZscsmBJvaJAtV7kaL2iZZtIm2O7sYzLVfL4LWvq5ijQr8
ghKqMPPi8hq6p0G6dJMe+5h0NbmTjrFjkYCtwFAuZ8BYp4quIzQMqNm8iC7txkDkyZ7N979cM8kX
Twu8k4Cu604fyltdSQF1iZCpkg8k2Hcn3ER2NH4KaGEPUGxc6d3ucCAWHWkNVhFq6nkVzdXGYo2h
k5ige1qU9EV0eF//r+fY2fGwlHTCSlL6mN3HodLAzqvOeaEZp8gWwhf/pg4+rv+xJG/9t06TB9KA
iQQT7oUXh5f5BYMfb/D6rnIZ+AiRRQJm7P1Yfz9odPXX119L6bnug/mPNtf1W2j8PFLPU7yWNEvO
PfLNhEyeo2baSdhJFIqNqIUVBKqBUVQPUuHanFe5334aXKx4gn7YiTqsekb7gEkLx2H01hJAUXYl
9r2lw/ucAZLzunOjj6T62DzL++8rlP9iFtPMZBnBDYHMnjs2o+dixFXVA9BAJgCTaF0z7UkyXkNp
GG8rlI9ScWQAqS3ITV2LGCmfoPVp8AAAMzgSudWjZAvgt0/tpCwPjXnTpw4IRjLTgrWpXkPYh2gL
Snq/ivvS5sbkttcgvnO7ce48/PH0Sgd39UjSj3eheK7NC9JxP1KgrLquShMwc0Y+WxKWFgyGy6Ms
RGferJaQz3/cnhvyW7U0nRRICrTkHVkZ5KhUcLkZqjY2UF6W6catQdBVq7UxODBKpJIoFdjFl9Vh
Gn7O43r2XnxPrTCa/egJck6Gq2zQVJmOsLH7yg+4KhibwiNB4ghaYUTZEm+MOPacq9m945XmMnbm
DR9OMtYFilEn9I966oBlHqYedit/BuBuANO1TOjX/EYthXVuhXHEta5Bpu5jXJ7Pdfyq9KsuWS4d
dIl/2+vRydAJaROwQbgZStAP8nsesmXyiXoQt1zRUoa8RDaY6hnYdkI/TsPObgiyzzZbHe+CkMXW
Y5WjIgyJSCRSHNNk+deP6XO+NzmZFPOFB3YAmIybbrMajXR5r93+6NWt8uoGcIx25RCrRfp9jr7s
Ujrq515okMGCCPSIykQzzBQ5jilfrnxQ6fh3BG2lI8ArXP+oPPK1CYjS705Tk9yf2hLDD/J4frHV
DJV+9muGdLdUyUBFayCAeXtj1QcOmDq7Jl6wBWWLqVQSp2Pn05anNwe3uWwkzenAl65qUx9NVZAS
gmJFv5zOpSEtEIWSp1jTn4DGXT1DsiE9L9uzfvnlxHAxV3zlFlOfy0doAJPBF6iGI9V8ipGKjidd
Hivd4lcT+FPS3TATcH8qlaYRX/Iol2kaeEOc+pZNJxzy/7KgEM7GCOh+HMtu3Jw9TCb+qDyaO4XR
iBOtMShwqh78FZpXjw0vmnZTjKEiKwFEjXdH/dwOqLMh0hbudg7Dw1tUZwgiqidRhiiWyyo849MJ
7JOlTft1GhuYJ4h2g0Jv39p7rBju+OqhriQWag2B3Dy94wGgAF7DcG28+2ufsu3Mmw6S9JYh7Y6u
ktLbPHAh2sll7ATKdhUX7WD2VBp62uFfuem7VahFEFT9OKfjqAsUyXQ0aU/cNcjFiaqDBSbXrOFS
8XHVyar2fSKAqznPoFbHxs3Nbo2/0eQ+J2BlEGR6JLeGXAZn1+Dh3zpXEJJOK4nyzxCoXImypraG
1TK8BwvHu4WwxamvZ60NwHQ1qX8HRYobQx8igtUQxBAsXwHrRQYyR64xNxr39cvZDKYfFkU93ubW
Y9Wrm9OJgI5J17j77pV5q6juq5a/8rwMp6xnBgep1bLLf3YIxmuqjPKhD5hnIpuwveMVNfIvBWuW
oXaFIDdxv9bw5JFuo8VnwOYvC7yEo06/lgq2o9OMXeDQ252EjmT38l3LPduTRXVwmlLWvaJfEGk5
dpogjYLrB37Vnga8+uam9aGjYIrMuvz+6HL6DiHd91YQ2omCczEZ0/zrsS+EUKgVUIRl3wRpsw7B
vEoSIj7RevaYHuZtPTecBk8Y1Gwne5b2CrlY3z3xKAQFWsxTPZEl1/SR5rgRTpBBNiFoWM1cjixM
YYm6yXTtmuVuPRpfRqW300vY3wHcHK+42SlZEzXdfjlB9EIHh/WTZE0f776ozfTX1fIeQkS8PGfv
uFzWjMx7BGYa7EsDsgIO7Bb/PECgF5n3lR0gyvS3qXpRZtjA6H0oWrLCCmp5p9FmgR/AuqMk1VnS
muJz2hIf+S4PUeDJObbF+LB9pIlpSMvSUuEj2qBLpxbpPckdtZFASMlFAIv/4feR80QJjktHqhbk
F8FV7nfHuBldr5e8w8aS96RrxPtT9bsjflVfZT6ddBR82mISuu5hYha5Hk6KAnVfwi2JSKqxhgZd
uoU/TIV3qMmKsSnpeaD9kTUnWYW3NfUU2HQOJXtzDXKoOQRFAjNYCfMw4yI7M0qRFCmCIMotMHj8
V54VLmPvowas3xS71ppNgzvwJ+z6fRhvb3tr1ewjd5f9ikCEyuG/vdFJSNL1HAV35maOP5ZnoA0c
O2Tv2hNsc3pfBu7du6SeNkHlR3h+/ypqM+417hR4cdEkrlo15ioinPhx2RVo1NuXlyRtru3axMDw
9aPLme/lH/hAYr7VFALv4lUNjKUjUslvmdAPHRVPpciggDzaWQ8GcTZogCncUudGy+AnOmlTMxBT
0ELrAzQ+mhf80RSVgXZetnDwQkmLQfKL/2egaxg9ouYouwYtkP48VqerW/awntf15PoYd8daAxe2
3NxetkYQWb6VqlNsFvhubyIrNhM86IRdJbblAHfZ2uFFZemoM4v7mSvxy47mxVYeaTekMUOQ6IsW
Cf7ZObuHFPUmIYYanwbn0URUoXlTYsPF0v16KkRAa5QqNq8ubS1JfuJMlmXTF3cAl/A7/d7HRG3r
D4k6x8L+eJHYDBac0eTlr8n1+hYVyNjLx9hQzfs+Bpx8xAU7wfgs2XpUZ2qi+6KCOCUqmNH+Hyu9
4X/Tistj9Enug7oHNFCaslbPeyp7dMZIgNqnCgbIcToMDs5egpPrSLLRjQB5mVV1PKOAHfQJHJ3E
mjJ6jIxKY2exA/PZdbt3bY1/fjHVuRB5+nW7pvGHipMPA9zetZOLCDak5bg9PZRUC0JDp9v9LDjq
Rd0HTdJnWVwqnSpJWqx8d+9PqeQe4j/75h1LBOjC50HdKSQqGTPLcUkXcvZcsMa5rZ2qjl/pY5sx
JNrlBwm2WoFgwGXX6WhoTdKQYTJ3ThI/AJTUR3MjQYaQhys9b32p10L9xItA+fFxCqAin3Sjq8f4
zkFv+B0IWrozfpqdfwxFQvs/He+pzP6qtvlTYT0e9tu9Z+ptG6hhixlD3E3G5qxRyF3ukM5YQWn1
3kC62Ojc0EHYTX6GIzW6tebUUSiegx7SpxVV+aIFb1NCDfNC05a4G63IyXk4682XctjSaeTtukMV
4sETeO3jyN1bofc5AppeqSv9mNYPIhYngAJ8WsNWKqLmSf00CgGoC8EVviKUj3YfnOuqX6K09tMa
684FXi65IoyrsvCJTtEK6SJxdX+2DkEsA1i/E9zgKVvAfN/9Cfyoeo5dvPSw7SsWpzU2a2iGqv18
K++xFoC1Vqp5ukAguP+EAy8h/uIVB/VR1eaJo4RJdymtEdG6rMsLF/WTAtzPEWCWjAoZaL0QxLHm
65VlDvwzhVy0YCz2YCWMDNipg0y0DNQxa6ITFhgHmm7LDhK1L/U2dDLPrdsrw/byXGolgF2xCFI5
8A58NCP5C09VD5pl36ioTh60MXophIvqlRJ/UcnNtqwQFzeFs4HA4IxJekH2vrr3seCn7LFs0NhL
haB8wegpkKMprQ7S4GGJFDMKoCNf5qmrenhN0v0TBPrm4A61RlTZUC6/4PGGrYqCS+JkYtmI7Yn9
QP7KVdzQxXA9bQB/c0hjQMheWMc5uIHSqPBsDx1NaZgtfbwEjLWr5vNqlFPeeCLui52nULZ3qUsZ
i9z6d+0mZWEXrcq2oQlvR/6c1roHpZsGkDbFeBJqfH+QOcgzN1Lc5Gawcu5rOiHxrxzINmlVCq6N
MRCBFVyxR7mo0jyzdQPEIwLor0vrOa1psYosWLQXhf1mnzDxmoUROEYWarXek/lMOMXRnFYRLAYJ
Lwo84Ifmo3xEuGkcgkbZbgTPaDrO54hz1zj9U2DRHgrZqESZxv6kMykNBGls9k0AnJ3ANe1M/b9d
9y70Il1C7Vmq+wdnbyNDU3nfZXcXv5fh2+BqZ/ehUA9c5F4ouBv55nLDZzAPLSGuH30dBhFrPeUu
qWUQ5s+PJ+mstHc194VKcx0H1tnasCM75rfBIN4P1RW3lwqK4wP7O+vdQ0eA2BzlQTINvrVg5EWD
B63lyISAaGpFoFz/2LacMZxbh8UtBORt7KogkOY6Rmsr8LHyEkVpxPrCarVn34qHOP4PwRclxt7U
MAZeT7P7FR2bPWT0xHiFhGCKkofphx7IYOYsYeo0ST0BruGLW3jBoZUOrKJ6J5HmXzayriR34Rv5
FfUfbxjr64fIMdOS4B5koN1QPO8sorV7kNIsJMIW7K/dzv3RZrYWapFGFp2fnVq6RWWTJHSxKx5d
ifhIp++HVVJD0DVsX+aCMQjieBS6TcKm0SIHSYRxDjBlK5eikX2dqE6gkuGWC51RHDC1WOm/RalI
SH7ynqA2pAW5vFbC3zG2Bw8tzadJntMzCXopAxzsXktbrSFKc/jlnJyfoMFZgyyaOIoSLQqgkfZv
WBeYfs/PClDG/pSfC09+wjmkdfnGTigppKwKlidZnJzYOxQxRPn3tl3Y7aO6W0UEAV6Kji2jph20
qWLKUflRNDigwY7BURj1bVcsZ+RNxatdyYxaO21yNRWzJ7jPTfqjJGDZvb1R93zVLT6g6NjF2wT9
XihqLoT5k3fasqdy0C47he9FjhjhXjlujLrlJVvKfLLWeVd0X5+CMXAJt/I5ZQ5QiE9+wef9TFvg
wC7xACgpuFCxDBbJdfgV71TZfY/mctQVY+MpibQ9HjbZoJXRMnVYjnfDP0zStbYbtHE3291M46bp
np+8dA8CCw0NfHSUtF3+fq/L5TFL+oHx5n4Eaql2+lcD7umZQ6eyc9QtIWEut0Sjgl6+oCW5bVOE
H4sEP1+s9Way/ybc4vsT5iFu8Q1fT6p2bmcSByDgo0+WesT4ypVq+wViZ7ohTf9mTAK02MTwQrJD
ZkbHf3gxT8ZNP2xcCnFk6xiI1RM+iHylil1q72H+7NkFo8DffEosdMCMVzj5E7XNNNSwyTXxYHSN
w6/KuU5XGnRho4Ag5wqTbac/0FbkkK5AkHkAW6zbQIaEHhE40ac4ZQaPtDo2hUXrGbm+jFLvrwN/
0GqriNHxfdiQmZSHmnzjk4UPjGfjkLodddQQKWpy6vxiy5HLGGt8PelrHDW9md3iVZXdHyfGE2au
uysWMiel3rcKSldjtxNcHQAGwKO5758gsxoBzzEM5eIZAi8AgwqOarlgnwnkpPTl36ktD9WwJ57Z
eekp4/M0uul1N1840QXeH5+ikvOLCtLRTPS2Uic2s7BxHvqaFgUhtdFIxwUpjQwsJlAPVIZNR+cx
C1su7Q0jDdh+8mS7mn5AeCRKlAw5VzO5nfIylAZhK03Hot/NPUenjNGFXZBMl6OnZZFkCaR6xKvh
nWzgCPtXJH6vhqsqlUFkiPJikTGd4iqLXWdVbTncaUgzpt3caHFR8Yft7iNCe6NMo6sY4XhHTtwf
Qp0Mq/vQFmXqAy7avS5sqOrZgVR3xQnZDm0yguXKRcAD69wsEpnzYcJhI43avhlBq+9EOeZjUdcx
bw3GveyuG0cY5PyBMKJA/+aMJ0UEQaM+0SUYK6KuaWygYTXDhV655nh/d7DwsqvLsG2Ebjy++Tt1
4jH6fpLfKF5DVv88/zqpvDgvjalYVkNGc0TJcyTAptTJynAPaLWXVhFxe9fPta5xpC7tMyyq1Pal
fUvMo4dz6PJi81dOlxPOnIebZP/W02k9CwUnyGpP6hPPCxLytdscVADem/+ViKoma74lPvd8hwP/
r55l4woWoTSHskdpB3VWP62ypq6YnDKm22HLk/EWrBXSobn0HTruDn7cGm2Xgw9iyIP1xYbuvZpq
ph3NZ3EJUmpmicJuVowoLpuNxiZxAlhio2V6+NC/5BmqePqAxNaux9Y9vSjPTrKEw/XaVsTtaBJ+
Ecv+JtH+m4C5kijpaYjVsreI6a3cyio/uFp0lutRmEBaKChGqBAsdRs12QH9OKepxvXDkwzJBEj2
HBaffdDPx6h0yJThQde9lJ+siKpRf3PDbiHtZyInPteSd0TXnVPJIia3gIg2yeeZuzwDDHqWIqGp
31HaMVPgk7O2QDCwRzCG/X2FqZVLFBk8QVzXVv3I1exunPGvzwQxx1Yog0PLHjw3eEM26Mk5nDJy
MZdHIWj/BaPW6d5xGr7QVUArDA12K92xv6glKAtM8Befwplw/MeXGKmp24yNx5O3pjbzbTRO7zKe
sC0ty+T5WeT7LNxa1j3ZYArb1xjtnxrJ34f/Xtgo6r9Eo+0ztabS1VzNDuBhDwBQvkB+8cYM4JOL
YjDaVoMEnCol+ueD8vgD3JKgvexqK519cSWppL4d/vb9rGC91JkRhAb+b7y50zTYxfbxkfI05Hf7
n3u9DWwOkxCN41ZL1qAuQHvM3tLolh/Q0K6HFEWTiWhHdjjS8eysClE86c7g3xmZAl+CzrDEFMpj
8d4AMtxwF9bkzl82w1PTfS3xr+CSrDITcdTc8G1kY8Z6B6j3iBZuSt9051qWakcrO5pu+cJl9Tkx
pecN62eeUtWGwkmux+F20MAhuhOCU+uNV+aF+UTH2Rz8Lwj525OYAj+5ogqGgyW2WtJoneu3P60V
HrUtrzZOk3DaGQZAmQZ9ytES0uCOA8yYR1Tf/LVfg38dhqpgAqyL/y+Ff9NBAGMq8aveRY5eRgtr
aRz55DS7tz/NbXx3F0oWBNN1ov3svpGKkJTy/P22qgU+iI5VEkBeR2DIARBJXXJ/00khfNQL9ENy
UsmcO7m17o9lNCkNLE1RNmWPNkSL7W0+qW2UTT/jPHZePoVhCNL8VqAJrHFT/YAO0yRjemCKOtYW
kMfrr4IQjeI5BxNmQCLsy/SqTjRmZ/oO6kLeOTurGFPkxcKqn43IL+IAWbu+NgPv8I67nbMKtEIO
ymuiqVJNN5gW6nyEwY8Pz1rXYD6k+gn/bmw1AoJgLKiT7K4hqygVHbnT2EfeVmkRm3/XqZ8rY4xF
jmHrvPU6rsOHs6r2vl9TVhCETgBr3rmfhJflPen7pWX44OmDmapXBTd4WA8FGmZKp+BCBYAvmzwO
LNdgP9alM1pMlw7rrgub7FyX5a0b7npyKSQztMox6c6YkMjU6mOJQjZoAuSoCr4+VBZm2c/dNp69
EErXI57IvU1/zvb5OIwkiDOOAnl415v+SNN15VAQv5a5Cpcj5FU7DmAsvqXhtwKOAxeiijPNL2nK
y1Xo8ShQeRWNquijHgjjsuvPICWsk6+TLmLpZks6+QTachYBzBXXyn9hX9KVieUBimlTu8dyduTT
w49Sm4v1w4UGTix8EXpesEyOAd//0mBaVhZLziux1OicURM7EY5VPafPLEndglEgxOlQdiZVjFiG
1IlWV/0/P3NflZQodsjaK6WfIN8JV2KGkzgWHJeDjhYmQWQyWhjC3R+gjUNLngi51LgN/9xTbAVQ
7NLESPr1CPrV2scmFy7thiccReC+guKwuCICO0qF0RvWanBTT+g4UVzt80vnx3Uf/9xsPE6ccMOg
t+4+M0u2vd8rCl1UlDTq9D4LQfTC6qCteNEeIe71P7KZl22b3XF1Oi89ApLr3/x4VANUDXUUwFp6
WtJlGB5RR2QcuDcZBLO6tvMHxRaGfQA5SVrgg38dd3tQtJSmumJQhBCLUQBWe7/rlfCfMrmqx1Gc
JQ81B2yBs83mK9TKVRAnvFHKCQMle5SJeI4OrjLdSdQV15riGSjb0TjUbiYtK5ZdvxK6K+8AcU8I
8qRwqHAonbuZj4Wk4uHW/PeYPToo1MJd6we3Noug8dYxzc5UbkMvWYW5/VFPOICXcQUXlOFWYk6S
5fISSdUfHR8aG5CzmjW/bv14B1m9O/m5ygAhhkN7VRgY2pfQRjC5tOfc6Q0kAw07yv7iQjdUVfTf
ZT38FKUiWWtAtPBr8OU6uifFmBXBARRf5Q4EwACsIk9s/WcD8UnHssWl4oLj8tcfYgAmUQ1L7mqo
E7kXnUGkNiTvoIQVjgsWlPo9jIZi3MqD+g2ooHSZMB5VlYpJFGQa9dP6DWaEFQ9tItHP9erL6C3s
ttLdRMAbMX5AoyjdTvgHNEggA66TPOSom9AFBmwRktl/BmMvStsnnOrhaFLdV94n1wZBjpYi01j+
jcz+ox2fz75CbmlDWw01wlGBiReYykCYTviqE6OQtLfWOEntwmo3FsquxkiHgdCmBh6X3CBWov8/
NBQvExzh8sjZQBqlrEbQktE7igD06uUpk7uDr8OEdesZ9NO+GOhN9IY5h6JPNpBGISuCbCWZr5FX
RWJsk7QjUghO2PAjMgOFpipDy9IJ4R0MhzW12qGlEYTb17bDvlkOkfEU5pj6pCJJj2YLOS2T5bPz
we3QmfzEBXDIwSqZtGzsSUQclcvqfM4BY+GndZ9pX3xZdY5sbaJYVYeNiHdn60IVM71T0A0bwX2j
pH895yIqYpCWOnaC64p1msZRpvUqjay7qQbiuVTvuvSuxA8YZADQ1HAauhbZIUS3mkndn6DldW5f
BktQW59t3EtdD8N5FoDD3WMBASRqjh6/8DHDEKJeug2QVGCTrQQhgWN6yaxTnhzKLL1YyJRnriWl
CSEmC/seCzpFRnwxXSpnlnXm6FA9dFGhP0yW0lTMCLSGwQ/PdlZ7l7dTQJ1DKjLk+985uphApPpx
YGRGAi/yws2625veI+GLqdSGj4bPtD5KoyOxWkWXvPZ9re5jfaFqrU6pLtuwb2hjUgwa+kSk/nyu
0eHiZL4jlqR+EZpxRFFcinCeVDsqfB/jhtTsdUeu6N7ogg8UjPNj+ePfBmjRE5U2IqL1r+J3f5JL
NEF8LYi6ozYSXRbLbcpqAhfF7VqWyyO90Hskq3DnhQBPQ8eaYG8ouA0YmDGO/Z2Hx6vh4M3IWpoW
W77d9vHtl/zX6zB3AVxH6oL4EgldTina+1ZWoAhIQA+ATS/Uv9tOAMVIPgFsCt4nBTAz3/uTI3rD
TPLVhyWlYQ5xedp5MsllzZsKomFJ8wAbSszxy1KuaHl6bpP0m8J8OfZELiJ2QgfvydSCR/FA6iiE
BvmK1vDf3t/dE2YAzIS3Y1orx8MtqnbVINob8oveU2kiu6lpvVUPqsz3JpKf5AltapIYGNG8uyqi
ax3gGjSVI/jPHBPSm2Spdhdv+OLqnT3LiU8DXmcnysX4idBsuj7aa96UIfhOs93r+PBBtSD6fBHP
rk02Vy04hZ2IrOChS78bJiLvjmXYhCA/JFb/fErPbHZqcPrBnPfFUoOmjizsNe1Vdgn3SuttNaPJ
VsSnewzgNVo7hJTNId/DSper5sQjAK1gPF9T7yHSaIMPP2VBROK4GQzF7avRxn1gtZDd2WgALMnA
3tsAVSy851XCNM/U54eJ54MWOEFmaNyvWQjWVxZfcQSQUqmhvLbPr6kUzghZNkI3CLMMjb0PxjlD
lBWlaluetal1GGptmgZX4dCM8UZek8VVrOfql3wLzTFrLkFdRoq5z4gOD9VE5dFIwEyYYaKX1PeR
tDSVaRdRLMv0wLFxSEuOHJkz5Y06kQOJnPnDiRGUNwxBu++9uxbUE/2uyTv2Q+rU7gdlR7LZZ38L
i5zqMn47gtWVAghBrXwQUTvsVTeGr6aHDTZUePkHCJWiU/y4dGiUCf3a37abb/1IlSezKdHGoV2B
hjZm1O8kOT5ifHMOCYEcG3u+Mifup0bMTCnkyC/rUD0l9mMeatcHWqOV4cGKSysIhXK7Cqct/5rJ
gacKW1mYzG8MYfxdW4xa2soVa2bY1LKTcLX/2iaVknpcdexoNB5pM8D1F005/YnAcxJ3tu7Ykq1R
mcIZs/PpPVAky1sjoddBAkOF1npsiUsvQzJvlLNLVxn+qDSFfd1f0sl/MyD9EYqsYq+LpdkzZtby
AxKxvaER05rOluuD0tpYTEes5P/7ONP6TdG9p10d3WvVVfnoN0dsJIyfuLkRYRVm345p7pn0oybG
Gxz2f2+BFGvt/CRucV/ddt6Lr65jcy3obMv2AhgeaAVn2b++ef6v/Q/Fed9RKhlH1vqUzOWDU85k
c/IyKo1kNwg7K79uViebXrKgxe5RIzPbRJ7THU5oiSPdqcl4yyBtjImPFcswEt/n+zR6t2cg2bSW
V+8R+n7XkXujxySVkA8JR0sHzeeV5IEgWxBGoXgQCC1SKgAMgXm5jcvz3tOa+RukMnDPLsvkxlp8
cgn5YgwoXy743SYm5N/ivhV8shf7GXGqYfClLU3LEg/lCNuOGJcJXFX6X5o85zWoO/VuiTBZNlZ6
BU2YR1d6bi87zFhq+8+1aNM86L0tX5WZVUozT5ABdb1lPbo6ZtDPwp3Ici5SQr2dTXFI8643zyQi
eIT021rKDX0YjXnX8vFv0gaCbSgCJkhqJ2gAO8TTR4A1drAnie32YGJT97umLCTgZT55j179a+hH
k/38lgGXWCHmiF+X1xSp3hZRGaTm08mBi10QF7lM4tXaP8a2GOw+mnTU2bXKFf9pPbXkUzMH2Q/e
jBID2CJig14k5SX61JQdGhm6XNIov4L0u87byi1cNCx91XqlKAtndDimuIFDqSMS6tcjsPX5nRg+
cWR7dw2ENMWFJazim+Ak/HoJVAE43YG3Dj4gpPh5bdWLEfzIuhRu/sweYgBcTSB4fqValtNw6Lnr
jyaPaO02VK5xeu05g6B+c35ckAxUrVyymZdqNMiWffRi27iHXP1oyhaJnZwQlq0FXOmUV75JWAfP
1AyRzxSC4arYmB+lK0JoKygyaSQuvnQxvCKkUBkEyZjBfw4retp7tdGtbBZPg2O0EndnMWTXYc42
afH2xPPaLx91uL5Iv7U2GZ+8NvtxVPu2IHdXbenV9+WprnNRQEUVgeSS4qjRdjFoQQzbpqh5wJlv
ssU/7Mn2KkkR1eLOeAIfCOxwAAv/XhgqU66e5PuY+TPdRdKyV/pL8hZMOKpTnvCHlAr6svYVorol
vN9dEX99eDNSjQGUZlFnO6u3E8lqDZFlgqtQY9eF8nexZQgetgo8BGOfDYG69jtZ+YPxsRsQK2Mf
2tWAsoky0OGxC6ZYfdYdu61/zM4B4tvg8oqEUzXqQVx96knh+YF5IyySASV2+cL4syP7CEyHcdKQ
YwDLddB+ZUF01NwSXRces0ivX0QDHODCygnaxtahoiTlBPCFIZz9aO2r6Ctn2KPrs9z8uxZahtPo
Nv9FqzlKPNxG9cRgg4zRa2gj1D0vwRicMFwjGAtnbjxoMZitwgafK1oPIuB0B3JMD/p+vwxPtm2a
nk4W/Hx8Lgb7nmz/LCSDP8J/6mrIQYXxRpmXBBzY5bMpCZ+ZUAxBVziirCGCptE1fxcJtPBrqyX/
defxsAzX6x6Aidssm669ouoTA/SoCDhW7vSAqts2i/LAHbQQyhAlWvT0sPCGuCGjFuqUxsoOCX+z
gduB4+y/gG6GEhPkvd/Su1eL4+M78fVUIg6Oaea8JWr1S2qQgkRlktYrUEndXQYaomeSdSuDqEyy
EyicP0yIeXoH2E1lk5xs8YwhesLdIPZAqgoJOdFz/Gna5wQdyYfgzn64m/pctQ60shHSobElpc0M
PcE6l+1K3faIOiZdykWzuNMhteLQHWJb7MZK5yqQ31BJq/Md0fOk4Egj821KZ4vzm7AVk7IJ0brn
fIJyZdHLQSwp/6nHHo8mEqKIQgthQdu1r528iAvI0yvjNHJ00LzzRSx3zdUCtHqChD5StXzBp3qP
HrD7LwVt5BsFFnADFjmt+dVFX0xY8sqJ4VMu/VGINJOXjxX4aD1rEabCe/8qWK2QUcvbX59oVMPi
g0PvOLUDHdmkaS847F7BQOi2FgLA90+FWxACR8yy3AhKTSt6mv8M9wrKBltX/OcbD+Lr1Rtebqrk
1LV+RXCqBe/EYGupdtb4PDuI06a66Xpl3ii+Xk7WBvp44qtL1eo8KW1Zd+Cxz4h/1gzY8PEAhrK6
oHGfkFYBzh+PKWJnVF56jZqTMjOx6Bd4PNV1s0UFTTR9WDYAK1bnvs/E/1i5GriSwiurnMybRIFG
9yWb4mEfrgqFOTtk4PEOiIYF0WCChAN+HVxj6cjjdJzT5J+oklpX10pKrLisgQyNk1S5U56Losjy
Ic1bT+mS4j3XCQS2CpkQVoCPSmD7gbje0NLoF/Jihhi3ySZCCDBcI2oqtKzKLDHoSsF3uW0lQAMw
DijGs1RDs668CvVlbaCeujtIUrwpTivn82JKh/LDf+dV6Au8ucifx4NqxjxaJw46huUR6/ThSDyR
sUw+8XYlIbTZ+Our5TYBJI4JlPgxXsKVVrIjfCJUsC17ikoKdqnWB2mOfjuAtqMF8oe3RtxPjV0/
hxIIMxBtsHK6z3h25Ut6Jgi/7o/XwfUBBz6JBvGjSueJM0E9dzb5qHHXtCjKdKyrn7aebJ6Rebg6
OQg0ADsHekJnebsBA4KSZkyreDukVTe4R8NJujV/iI0iIGJKEwXBQxAJEV8gjAzjpI7m6hLyxlOe
29ZE0mbDCJqt7tye+ersf5vmzgH+MTShyF7/n/9O3RwztmUlE+imjjw/nflA1nzshjBI3oLrDkH0
jDygvL5+2+JKwU/g/lf9u5tyqdybBwI6ewfXAHx5vH1yuSr5D9mby0atMxhJK1RuTBbjBGhTfhwk
A7x47myuzpBFYUw1HRAZ8CtU7WdpnjxDSYy239p4kwoc78DAaJY0Y4vdO3AjUyCe/C4Pl2337gfM
pyJhjGDtyMmpZpkDNof4uN22lNVCYhsy4LbY3DRo6mDrZ99uLS/R6Ce+8TShbWi4j768MtVVp8B6
RKWMwDyDrIIw6fkIVDndnADQm6aouaqVX3iR8/Si+A+6Y+VHf9HtS1jd6FigFfn6z6JsQK+Rdubm
hmZH8dhIF7D+i8HFXq8sjPEq2MNIdum2pLD4eaT6wJYFLr42+9+efpSXK+5RbnHebCnlC7U1Sys+
tS5NzV4q6vWDDEJ8eIUj91qb+Ftwdm4v/4SS5vN+eywKJ71D1QLWdN6ZiQ7YT1VQgIB4xAhMeOAt
aeDQnPwo1/LBq3hNKmfvwi8Oq4F99/aEYlWF3FzhKWSM8Db9a+X0WkvKiDyIwyAhQ+h9aUv4IHdP
gGPhjtdrQtCkRghwdQ3Ft/DgjLAowtZor2gLJzmxsHgYjTVclhR7SFW6xG8C97t7FMG8aZN/B/fp
E/bWvYpZ7fAIqXBgGWTLvqrBlrWQuxAokqmyktMCI56BgK4c1oen5PgB0yh8w8QttsdOxZSvCYwh
rHzjtnlZQUtXCCuVTMg7u9a2hS9ZA0FBHSg5Jvc613EK14WBgpEE4mkZFNqSdcKmsO6PoqAGIjWJ
wmPIT46Z+1eMf/gG/62FjjRIY9Bu3G4GHirrsd01VwpZsrEpj9PwPdc+v2gp81rk4IQHB65AbqV6
aD6jbIC5DbFe+ppHFaPa05oW6yufWMCiNebfa5mftGLbl/mDguKqToNoNa66eiSgtKCaHSsa5FqK
BzorIy+afOVPLpNrZchqXQyhfFw52uDGNNrZyvcasQLevNUR71JkEUcC2g4Rrvr87ivVEZFx0iyA
fOAdsgPxwphw1pHMbo4MlCEkYgXg9SDQeSs/uAqNRBYOaiikfhRF7xAnCq7OLSqEgLmdzQor3QUI
LLxOH6yv0aePpVMrQsG1ZxD8VpP8R8CLQ+cnbrmLWXzg9DYn9TWh2vqxYIeIfDC4IbqV1fTgiF2u
cafWasuHk20qtqdfdTP8Fd5Rn9DzeytanOvGJLAdDzd30RlL8oGFYm5vF1jkAbSQIkh/yV+Qt/3T
J/bIxEHe4Kgb+WmNrI/LkOLG+w+5RxXNzy6lKioT2z/DYKucFLxOREJ7h6o9IYB9G4luZmkYz7ce
s0VBAlBJf0YK3xWHZJXsD0BpVceR8f9wiUKCXqnzBoz4YjQg5BTe9uooRMLBiNdaW3XpfDYSmojV
yoIXa8ldbkyozEavfDGNnAceJieN8YnjNL+NrMBimEgjkMPYrl2t5OxUfc9uh+LEaATD6mxi5ZOy
FMNHJoAe3WJMsm0QB6ryXENc6A57duyFf8ZpUwdszy5RzshhtXQwaHy5hWcFL1N5bxMPAtRW7K2J
d4fhJHWLIjAfrzZSjcxxUmi8HtDUbuupqJfYTGPFYxKWQ99YvwmQG8Ykurmncqy74oZPyyEk8xC2
Hl3EX04d7UX5RyjxtaREsu9OKgxmN6iTGtcVAKxAeFe9O10pj5d/Y4g9W6EYYEgpPImmzkNknHKj
PSxYTKcB2XE/2eJ+EVf3zHlGSxeAOfkqz0rlsK27TWhUyx7uy09QtVVugiRfPxMjXaLYzMLhaRsi
b+tNSgu1SBlXDLitupRXloyKMKUa8qrlOSwpk4Ljr9jltmRMv45cEUALIOWyz89zEUPHtuKj1Ng5
YpH2R4aiwIb5vQ3WR3cggua8C8UmwqIw/OY/fan3u/fJVK9Ei/hZrAHXY9sx6/16iFOrmVkZMvuL
7FYKh4VhfKCk3y+CSTa5OMxkdwQx2Bzcos3iJ0VFnU6r27tz+1sWtuXB1SLhbQE91XnIG6/5h18C
/kp8leSDxSufDUd5Dye1iPxI89oBqp/rYFhbIfLLu/4Hdwp9GDNBRw+NzOyruJkGAIFrOdSPZE8P
rRkjxMueTpMlqS4D3Jh8Qg/YrF603tXzOAZaX83ZkqqwF9KJV+e+g2S+wi5ferjmppYAFp8EZd5w
8s+2D7ufJzP7vn7ZsKpwvudhCsPCls1A5ukDkAE3ap6y8ujtSq+8M+iLrlA8hQi/264SEt4cWkex
cxnqI62dpsCVEdYJJH4YyHD1jcG0hj+IeNKskT+YJ5CEYzWqk8TGUFX2lc/M2xboRHWj+vqriOLt
Q2OJaWTxnOad6ZKn9hIpTr52q32WFl0uOt6TqUxxoFwI3qvcojaLcltbloRfBBh5CscFR887ewm2
xM1+Bp1RCdQTL3kCr9Vw0jkjkBvUUa4R5zqP1JzyToejnHi29RfyLhKEVClhnUVYl03Pj4oo1FcH
yrFb4IRghvLoMg68ihYqi2OvwEB56O7tkF89/lZoN7ftrscLKFl1uhtEvPBzLv3PVIa2tGWF5Rah
TSEjKpAKXJFEUQCoP354Ra95t6luGV5Yk2jFyXhXrqtowRcIl2HTsBw2rbYRAROVADKFrDK0kBCC
QA1GN8eFI47b26pCHlX7YvSBjTM63Sg8x55UkkrAYnphSPqjMbmEuUcc83KBT/Yxoxn7rZeJv6nv
9tVBG2nMEmC/DIx1OncP68nhPTEFm2xRQ2c+dow/ifCujIu0FtOJaXXW4kiLy4ZmPLGmTxwyw0qv
0AEr4/dn9HbNzfE2CAGSudzKhMuMqMjMrhhJdMmxDF3/nxok9xqceiGLuvLLbOC8+fsos2SdCLCi
g7Ah0AcojUuBI2M3s2Xxb1aYDdzY2kGyIRai+pct/UuDPcakOVNHtDILYzH/8vLP4x2pBH6LBBB4
C1bauC5YVGvDGOUC1/fZCJffZENH53tDwi6+htkeribAQP9PR6jKemso0hS2Zg/U+a1f4RqBUEwk
miKBPm5HfzOzjPligcX6NXqbAkTuCkB1iJIzZogLNNlfjwKftUFdQD79YOJVqP77IpN08wKliKAt
R1QSoGbE7Hxs4bg7Q2Q5hEd3zL3iRDq58XXcg0mPLvlvdeoNcbZoiXhMw6R1EYkuY3g2zXq8x5A4
y+9TbGabaIZvrJ6zLTzIhvCZk3EJElkEq5B90DLFxdq6dhJEszr4gSciGj5rpCFlDIHuqzTiY5dL
pFfvjQNYI5L514YthhNf+TYB12W9mCkI7pgV5oXhidMd7ahJGX8Fl1A+mSQmuD7y1Z/xvknBBAMD
JpTurVsZeFu3CBpt6sPBS6dhz4JhxhfaG8MvokYjdtFRlRRAT7aA/bgr2jRQEu9A41+15EC2Pqhd
AfenpuxzHKT408eK01znW5SoSAiqPp2UJNTsl25TdZha6XZuG8t/82L7hRyVGV7MD+YETwwg2glR
4H+ju4E6jHiunATL5LgaCIFCa3eantI+azitSWLghAHPxunRrnfL3n4WuDfr7DWV7NsuAOgRAgcb
eDwZCbXImZWxYgefRmdjdCb95MxkwB3xRT8KComgZsPASNbjMc/xTht+9c8JtKgpbX4LEeC7RWMh
LIsjvPSBb0WD5Ng1v3bbCrKeC69cK5Lcpfe02+z/OYnIcTW2oEflKae0Ukov5PDkVXvx5UEHl3ZF
aokwSUF7kK5L3b3W0q66groebxuAILLf4EjM4AmU+JtinxFnST9xo495WkUO86MusJNo5JuNSByr
rLSXlh0Z50uP6xL5wiqXAj7mRsdTjv/cIfGIYIvVWxQyzXtYIGapXRQ/KCPW6XSq9qWDJQDpkCIe
GMCHCxmrmfioja9HsOjnYcwIBxlTRDHZ23hITkcGTxAeIqZZVi6MwB3NKvzlAO6heJ3q9FmNGMDB
nZA0JYzvSQOyHUVZxOojzrgW8avQFhr3n/mbRmFjD9cetdfsTwHPMjPymCb/vOLBbGIX0VIOI086
UOJn/rpAu7N8ApnFe41XxthK2GBGxR7OD9lC4dlaoveqe6av/pG8A3LOIkixR5ynhnwkrpUaeXjt
NS+KEI5ZYaZZ0p/lZxb9kYnWoqN8iOB0tamespGNg72zQOgmDJOjwo3BAg9BDJKoBoE2oIcBNMfQ
QHt0KigaFKoGfPE2GkJ7SIw0DUEGajMBb472ZNRZdO83RUH8X4JBTQ6c5+F19/slSG6edXU8Qseu
ZUSO/qYAk4qwF4jXIdjy/BOxT+jpHdlvdsrSgkEjdIOsdaMa2EGywvrWNjK9+PtkJK2D6D5sdjh5
fK/iJBPmOY5cFtMmqcxhZDYsVkjiHqBBQeUBjY339eyit675x5yh/iMRORg2YIgeogOJoFW8orWd
dcb4u9lOGhIufGHHP2mvXzk/frLRNOYYPxF+LAY///HxDRnwjYWP0wQlMTS9Use79JiDN/UoZLqm
j5D0QHSmiZYLSDDjye80IVh79ZaUiOQlIIo1KzJR3m/8RMuvUE3tmWlcjN2vpu+QBZR+ML78H/bb
tWORbMK4cxduAQSOGhczHvwWLcWgMQT6sDiLS9frvPh+a+uycQ6jTBKI+XomkDj9ydWWjJYuYW+0
/61srih6CcE4iB+XoKVkpzO8hlWNToH2C4rO7c3su4aINaAk45XnN1GA5yD949gF9+EG3Ox9816s
sETurfNgLpEk+Qk7O0pd7eyQZB2cymn3gNXv5A8JUTmyhQU36dgf9Rjvel8i1pmm6Q6V9IjImhJ0
chMt1/Slwm6rb96Y8Go9fxu+oB3pkURW4zQUe9DoH895fCgv0Gqitm60f9GZGAomuFMsmvwiI2P0
ci3yiDpAaa2RzwpZmYyD/BrZ0lzgxU8pSCTe62iXP9LTDMCkewEEbW4F1h6fgRNK5g2p/SQHn0TA
TfjMwKYtUe2ybo+B2jBSTF3EfMuf/jiDor2OHhFrfgPZLQ7KTdUDfvNBTH8o8kKC62TUh2u+oFKd
P5Ct4/TcJjTEJ0p4RRQUdxc+rJlP8BpSktNq/2e0nzx+VH27S6k3MzifBoxjnZGBgKOeouRILLR8
oN3xA2GAC9JjRy5fJeugHkJYI2PWerpQMMxsqHByVTmpcv4STZ84CNLsoZhF6IYLbH6Fn6rRazke
dAlgbd/sjMnXe05oVUlF0wqWgMLlM7ydTw8ZNtSIyXyF1LV2iH02sY39BJS7Gr3iz0Xgxe6kAix/
uGSKDzjv1qPKeCGknTmj+RhR0rev2JDsUfzCioOxqIM7AgY5JGZhZb55ucJ1x4yvc+YeLzv0l0A4
RaaOaFGzTcnKpQ9awTDiAnHFxhNRRmqNCNXHsma2jofj1Ledy7WnG4fUb7ORWhEtIdlGLhlwwb88
5B8ndFQwPiLFS1lVI5GSsaL6jEAL1MXVgOh6Vi+jRNM48iHNTI5J3j4U7Ek828kC0vt4bZaUy9h6
2O/mCy2Edvc7PXdL/xzKVs5nD1dlfvaNpVN0b/+xRXcd0Oz87C7lS9oH2wapzxmBSiUu8S/djmVe
T5IvDXg0bneb2vigWmrwoUF/KISH7NbpbV0AxRpuOO8UeUbsa446zKRJ+8rzQkiNMfPU6rRn5ZFV
wWfKTghUA9/JUd38n5IjNmN41p8FtpUOc6SWZikwu56GwQRx2C2XY8MJq7xuc4qowufswODsWCZD
oEOtsPWAqEwxbkm+XhM7z5j1h3fUCoYGKpI+MLojlkdC61z7CSLc6rD+jQhtfH7am3EHe1cD1cvE
oD/6lNAEfxc7wuf8OdZ+CqbdFUCFPQZC0gydi7NMw8ShZxTcvauVk7wkZvUdyIqKhe4xiMMW9nCc
JoIhhHrEXEU1LfljVlK7wmLTQE4q2bGVGDgvkSO7rOtuQFK9GD9lL0J5CUvucjo59/iM5znKv89/
QEFhNOb17TFA6qqjafOs8vLJ2iRMA/+PVNqRBmXGDsP8z6DVW0HcVQcbGYrIKGPoAG0h9B/F3QQj
tK/Ji79N4SmMQvd2C9OHPoxGUCtABzMUUfNFrB5bnXRHPOUQ+8+I033awZ7KTPXHHgqXllID+lrv
gh0ia7VFviTKFW7+ESvNwXqer1UThEtz9mgIE/QhJXHPy1V42JOmTa3yUZHZ1SHMYtWOGFN/gGY6
p3q+iroJcUX6AJtdu3nYcTj/Qbi9451IQdxH63XeXiCcU2sNq5T++o5hFws6SsvQttVlBwMj6Grr
Fh7x+k1lQsfvpjp2sxSguREzz8JuLCFTVZwMZ+Pnx5DhTB3FfxNeVB/3uaNzEpqJdgUtyf+gMDLn
1Tu8HLZBd833hi5LsgcL8DMQx0wx/VXzD7XCsuZY28Uku66nL5CxMBhwQIoEsrvjRFLDYsnpTua+
iG7l9T4xveoABf9OS7neabktqWjSDsLii/8G2dg79OTnf+1PbIJQ/1JySX7xqh+oK+R/EahDvTHZ
JXkvq/4VZzWX6j1xf/pPe+ysH7WwoGpta4H7XJTXVvE1MT28VzRyXAP4ViWXze+t08DVcI3mb4Tm
2+YFogTupuSd8yWzfbwB6GDXJv3Ax50KXvwrg0RB681fSY7R691MO9CAGVEaOzOGrp6lmu0p2F0M
tIcDdzCw4Sdb7f7qc69lgA+GRc0TPGK6PKOAPseKXz4uUWQ0zckHWCogyHg18EEM4KTITtc4omma
LXctF4RLsSZmEZb6UFtdG8YEus/U4qyrjiqgM74lf+JSYGreZ77Y/aO6txA/8ZVguMGPzxYCwDoI
K/wbDkIUKI8PkQC8ZUAx8wvkVLOq8RNevDezf3JmJhEHEEMbUoH9bID+BylNjjLX1XSD62lm4MUm
BLKgh277NCw+tsE+XRMEMEGp5n1ADkAZ3EKmycYk+lZSXGGkVk/Ujk4xdL0oRwaHvqFjB2+s6rpH
ByfFScJEshZD8K0I+vYVfNs/312sWw1yR1MdCNWYHmj4wkzd3fGNDq8rbnjOjlEqhuvbR4uMo7rc
nGBnTLk5kOxUJozdRRorZwLxDGwcXGFoRXhwqeS7v93tpzAeaccf08TIR1suoa9l/n7dDbhAts1g
hU71lUEbrXMyAH7q3wT3fZAS8YMLT3Q1+QeoUXYgFMRfHsBdBXYieyxLiW3trfDbvVyHjHalN4pr
94mNgQFoDiWvnHjo4+kn+0YFBIUpRN3V+2cX4gNSYgMHfWBvegZje75iO1fEQWKlqjp/Ya/WN4yP
Q3BDbmujX+yvmgwbB1PP7ss0loO9iocoa7l+hEbYWnqUzEia6Qrw4QbMx9PISKoZTeDzUnMcomFw
eTAogMwnzFHQUrUq6TDaj0b1+VkCjRRWOJFHv57DPDGT6BqKeoyMfxx0pLtF6sQ4Oq9NzCdF41ge
HVeRnatcAGPhdmhiOAAf+k8PRzUf8+Qajd3NxT47UV240J5r8Xc/Az7Ww1WpP9FU7mF1JFH9VVGP
EI6B0VcNj9paGGgL2FNALoYVMFPLjNMc9pUnzpieKg/SPVEY6wAay5TOVzN7kVjeU0J2Kij8nxr4
auMezrEdxckrUY/W91QSrXq0oHM2H9AZqNJEoKnVD3hLSPzLs0TAdiWoQopep3UwIgJw4+E9kbgG
ZLk490qz2vaKKqjuqx2PVxhTPZYvQZoBSsM0qaC7+JmcqYsGaXfc42SyEwbDYmMDZYGISBYghgm5
pibGpXYdPL3TD4ex0QsNixgs/RU5SgOmTN7RslFjKZITUHdBAvgP2NdexHCdJmRy1So26kEFoDbk
PeFcUxvsZ9hR1lX2IXv41sUPcaJID3llJ4i9H5WLIn8Hy4IABHxWzYmJQzHtkS6eXS8BVWIXSUNl
RLnTiEff3yZDGh9xP90NwEHW+g2uvgz2YMKmTUc/ksgezx2PfM+WTKJzei1Tj61ynXJbNRMu2m9Y
B+s1TnX2zAoztlPiYz+GrPSYHH98l0e2IVzFfYCOmqV7oZ92Z7PUDFxcGYXAChsakmiPccD+B0TV
X7uDIlQfwRE7ufHodLCb70EtMh85SBY3krJ8HyR6fbmTro6s5xpFXeuTqyEpNj1oFGWT6XTBJuub
nKYJMJDbBPUqF3b9y8slZJjnwr6A4nFUj20mi3z71y5eGyMzOGTWNlTHYgpKSky4hKjU4TjKfU8E
G1NPy9sc1MLMyEY1DEeYIgieFMyyLZsXT4H9OTvqWiA59YUZG1dolA5Brz7KYMmsgpHLf+U6CdX7
K9EvjxXnGn20H5W4B9t2m/k1KkfAROKeg3uj3aRo3Ljc7Q8XiVwcdrC6EhBDzAvLs8PTRlPtlXQb
6xXm9QvyDgO9TWcgRS6n78rAkndBnnGEFpk3qvjMINwz1AsYNyh8tlNEf1CTXfsDN5yGSeAsOuB7
ZPZowGj3GSXQxKvZBwTUTcsbS7la6sHEIY6UM8UBoTZnOuY5nbMOJT0Cl6lcPnpy7dMl+R3uCg8X
U5UBMpO0wmKJ83VAjijic+QQDuUy8zxACSItOf6vPdKzVu7MebyB9qnfrZL/XlwIJWoN099JAvV+
otlnUyZxwpmVnU0LBoZXTbhE5phodMR+NX4FQfP+TzkwR6k7gXZKKET/L7t3+0/BJ9aIZR/2pIRr
QaPtrc3kCWKZRfR8SVNeJs6LsOsLg/4XkQIrT6wo9BdVoEv0aalnNFukLA3jfX3EMI73+jyg+gxJ
GfxoB4Z+ODLvS66rNnf3wNspRAnzmL9LTE3EG4SFIePLRWltX2khVD8VPXUGkoBgOEFFqiIzbmvg
G5jvNX4jwytxCGlZ/DUFofdHSCEnvhoRWSMAoWaotDTVCPGe1UB6wOM0sGqYSAJ8yqWvDuAheNs4
hz+peSZMgIFcFqiClmEadyOF+Ob4yx+GB3EWhaxJJ0TC/B8YCRYY27he16vgBwrjbCKHd2SSYswM
pn5/A1HYjpzGHtuEggrYdTg+KVm3bR58jA7Pks8CYFlhMt2M7VJXRyFI2MUBRwpcfE7RKPo59cp+
pCm1d8MI0n6kRYDnSkDYTQ+q1sqrfghANwt/Td2MNiB8AWM2oQP0Q8iWqxCq4Jj6PdoIf5dy8sV2
bq6VcWhwNYPsahrMKKS7sN+51L0TqiI3G3m5G9xCdxNmS5MVlOVGd514cfSByhAJ01qUAn+bXwL8
TqcVILwy7fOTYsjGl9z7H0qOC4e4Y2oKnSl6K4QUQDPkW1es5yWXPGTv1zeMoqQLKOYFH977i7+t
4VWTE1B/Wm7s4i0iinqKEm8v0P93M5aAF3ar88r+51uHRH48rzKyIGDR9wwr7xbMMLPNHQ2eIrVo
d3tMDJT3OIg7QyaoFGkgfb7+FZSDPXrvHVzS77/CKM3oh3KJkhBZlh1GSrr0eLg71nJrfL1orQFf
DPTGl5+yii2T9hyJqwAzWQ9x7u/t2FCP7VC5v03c4UYe/ZgFx9lbFtN6rdvJGAPOTXyJkthnzfI8
BT9LuUhluA7X/ZNK5G/cSdEiHxUTDuDehU5AnsqSKusHskyuwBodpzSg32HfIdBtrkLHEaaL+ZpP
P6Ia2Kbhcz1wv7qBa8ruqBTO8bp54+h9uMmV7prauQY+dzf2okL+bJBBt2bdLkMpF9R3OVc1k3sf
R5me55+j3rJslCTdekDcHoM2HmRDSQb6weyPjKOM4m9aMVv2gYxM+Z60XIbsiBtEPM9d9Dpoqjpx
QdXs/W/Hk7hKprOmZ1IxTjKf9sLwQcfbq93anWuP25cXcPqmZuVDWi36tiuS7CRjxCK/buHEtt2k
GBZCTwV9ooeRPNhNmQR/wQa3EgsxoMBO7PeMf2k4p+19NDI0tzR7FwuGRK+qpFvhhXfvxe/QGMdZ
+d9sBSN7OLpHTAxVYIx1mvg46nnLIcYtb32OZr/HoVVmgFyVSCvjC6l3V8hqCnm7Z4ypZdGDNQRT
3jPxwiJep1PlRLUXDcfJaLyJPkUgd+R+C1FNw1hQtEJZ0txaQldSFZEUFIDeo8Bv9EGkyPSatJKx
IUBpdWLL9ZUB8miCaBEQgKrAgzHkr1a8fnlTD685gx7WYWwoC22hdi4+HVcUpSdUW1loSCM6yvO7
qJ0TK3GFFMRgWmrEAA6GSDDMOGU6qtG/LFFDY/2+CmS75KrP4+Yrv7otN7+ymoq2sDYaev34dUQB
5eCV5KNNyw+wmDnNUmfhs3rRezqOI/2Y7PV20Nq4anhNWdmhRWMB5Prdl5yGEqo7unCkAmRDKxyK
vqbhArEUiYgiiBrbkfSt5GHdDhfog8qYb3V9vKTtA+aD6VFIcJ215yowLQX0ivSzssTLUBNfNYMG
gq/8VLZI3qP6AKADYLTPCh1UDHPNaCTNT7ymIwya5ml85529to2NnQ1AFt8p3SXQ2JQPt0T3DrYf
u9Db/qAuvne25F9161ApKcTv6RjTuaFacg6v2a5FVJoKfzrEOqSpCB4/4/dIrQU1/LPgEAVtj/Zw
6p9T9IeRJwqktNNqkEy3iP7oIcFjbiAdtROz26AsGwH3Er1JWTE5HfkNhklD6DlURFkjnhKny9uU
PGEo0i8SlQCIJrhDnzWzpL7OsoA3fCwrDTSkb8D2fC0IQP1sKPzRIsgpc+afh4MpwbzftZ3Ey0n/
trKPiG8/AY8aMb9ycMJf/mEX+b5enuQvrb7Fst2+XV2DNLSZEjT4pBbPlFojMQObc7S1k+4WW9R0
zjhz1n+KRXpS/hoWc2UgfcDmnsQRtzfeJcykIqUenSxP+qq74EJaLf37QN+e6e+rBe0COk8ZjplG
tYnsb/fYAB/nHNVDop9aDG7oSK70BlbobY4qRo3okNiacMET46j6uB3rRYkHw8ucjxrCKH7+fwCD
+I2dEPvGahgyM819TrDrXRTXsM677Lz4EAMVCA/SBmVg30ZTPF784FOM4uSz7hn3ei8gt6QIOoVi
GN4u5hkl0yckBXOPzFy3a4pji7vCmjsHoTPsWc7tn3v1NGlgiI0BXEjVtjigwnHH6XHWujD2r46s
QDVREfrBZ2AzC4HrHioVfuLSRbNq4dnoGsUVPXzGKT1x/PriUiEcBPxA0ygciEklsYRnnJWATffj
jZqFafLAOePM2u0wQmpu6pdt/lP3q6iUiMeQZHTQztlnM23C/A4gu+bmI2qO7pDv5g8LSb/43hKB
u3QmHsxbfg3zcAUdYD1JzkB3vGLukDAFktUsx9Ibve3/jn0TqcbcI5CF4/zbm3XGJVLSaxR0XYwg
x5bjVW5qOPbi9XN0s2kNG0tawvGMECmgq+qQI1PgULbAWka3hyIku/ljEQNzYJdZoMlde5Thhg0t
wOFEsuaQootoLnBAoBFxmFimeAdb7NJLOloWb5tCnG/1ZNmVExoz6mzMT49lI+bWOibQVX7FDPLB
TNTJ8LhXjLvbyFJPDRh7v3Rba3NHoyaKf/3ex7SKl/TcMmEh0H87DsMwYeArUQKuIWlEy1En4pGX
ptlM2rs2kNo1IROBgQsMfuDWpCXFBlMXPAkEkNAMrlr0kM5Kb2sKpbYK7nmkRNRLm2+52EBECvzm
O2glzkHdQmkjZTC2KW8EpwLHaub/BG09iBPHRRJ+1WRGGR7So3Ojcin9fqKLpk725lEuJxOKppxp
spj0TUAcCzsAfaQMczumf36fWIQIZhPN0/FMYuf5cQTmS1oJpA0P5zRlmonv8vk4wwHgMeJsMKf/
IsVHOzebFCsUly8K89bkT0SJcGiz/aGEpdVcteeUGUrUgmfn3/RClPknm6D6yUqeroaPWeUS5BVJ
90JDnJ/5U0xFHZnbpt15PKtt1SuQHBrGHWV+cJnrH31sXEZxtghMjMN+IoGOZ2LhTvtylDY7MOr3
OZQM08EdALSkH3K2FoFh9Ifaizfo0dxQ1djLxuN9JBunLAx2WlaaJlYKehHgxopm5asi5wrm0eUY
Kx5L0JqO3M/UMDukZmk1SJUUdoFSLzCk5wgrF3ioxsg7nUwoNTNzMJSuJfZR96ffJ8I0fqr2KBmY
D4LITE7V4buXrEY5aBKcHhuLOfVC8ieZZZoyJoHLSZBNP7WF6xSKG7SN2wn4Bxoevbohqdcv20zu
yE2k/Y3TC+djcI5idGQw6BwxjaHOm7P4yjXVNhawI5vbeFFrb2h1Hzf+bBP5b1JD/Gf8cbMY5WDc
X8pDL1Td7JTrzXGk4+VU7VLYL9vOljWRS3siC6GglDPszq/oixXYP3H0e4hHdJFdi3xK120eGSc0
R25lCUokqmd46Tym8XDqPxJmI7iQgHUbhJy9un636/D+FGTyYAvAHuJ3+XPW6WXksZRl1RltVoxz
kQ9RoOi9gdyU2/9/2ZOxuMsilFM85gKYVuOrl1vkOSpKyZ8FspAntKJbhulOzeYrvselghSCT3iX
RyuydDydoM9Fue4CdFXbMdxBz+T1ZDZ13VI/3MNyO+2VCd+ltjo3QjLuxsp8tknsKiVLWjfWvEq2
sdOWSarfNXM15szg3nfGqHjrvNmpDE1kFc2LeTghzAxRdK9tIU8h+5tJjDJkCbB7Qs5b7qcC8JKQ
NRJ1ggr/OSXi1EvEyYd1f+WYiUVHCQS/mn6b6SzeXM9wYKUq7OBFKI9cZKl894fgyBDmeofsgRMh
lMrxqXxYLMn88mFv321fUr9Gp5UcJtvaB2jvZidExpaUEmdFCAKlHhgQhJqVGbIUryfH6Z30CNPL
ralTzRfd6ugmDzAyGvh1mgqnQBba8cIEmv+1HISIGWmn3g5s2oh9mfY2IqInWfQUM9fhYRMTwyLd
ppYutWBd/XhLafC5oLGW6uQsk5b9Z9nELpHcDbWSKsfI9XSgDoxTuM3EHNtu98b/oNGzo7LyrNnd
Ly3/IooMIjpEkrfDU1f49oYdzjMwv/1dZe/Uum/8QqwBtVwhBN08AHsfeO6zwjJgyEv7dBDXUQkM
1GtLjyS+bqHgO4XK9KU7Kxly+DGzIZXfs11r/qpM5R/lJUKIIzejpInAgtZDAB39U+rhD0LRJD31
cHFF8Tzh652d6NwQ1iK1bViYf10X4gS6ayk1zddQBgMndxHX8DUwgWhuVceCnl/uPVJ1x910J575
dTtIH13veZpnf7qcW8f4Kn45TTeiNBAXmP3Kz5+U9gy1MLdnb/FmBphvczHr+8mvkrEmDWoiQpvm
Y88O7ZeyWNbX6sjAbFSC8JrOEYpLcv+sy19Z0Q+AdgOFeBV1Vrg+EHM/XW7eyuNJ4jeQT2UtaiKB
BY4UPGrsMT1phHY3IARv/nN68YOWe3R155SSFYGm5/vu08gkXsJ8RyJP1BgQWVqT2RQLnlh+F52I
21mMFoJ5qiNsBF6RGSQEQ87y9j3+gP0V3EMvhMvTaC7968Rz5phqjN2GCBTU12bHUYAHsr+T0Ib0
c+MA4Rkk5xMBU/jeT9z226RYXdTBcVEcJ7SHuUt2+8bZCWbh1/KECvoEL2cpo6JM2uPDGvlqiNF9
2QIPMW02u09RVTOr9H2WpZAt7esPCpIDl4MQNpLFrXyllNIjfw7q+/Y40wKgl1PIXWRCaGb6muNh
bd86vq9j/oRfw/f2lPCNHBtBNZUdx/E4tBsCLzlMQ7enPwIzqSTa75plz0xeD0B58u6oEZRRx5yh
VMyQTIY7fn39EjtOI42Arzzv7EcOxzH4BazT0ydHymdNM0bAHzPyAH3vIpCvhC6FcIcKTvRLt6mJ
SmMLDM8vcx/5rO24ODpkJ2cMqmTg7OsVrgW+lrZhrRn/iv4+jXGKFJBmYhRf5IE0vySz7aPlWJPs
Lndej/JxMHsIMU1ZMTSyYRRkvrQuNfsZ7DvlDQhYPF7MDoY76oFurdDcIVpOkmFewe7Tr7zHDAA9
2i/OdCoS4PYWuRoSsx3UgCtAPxgk9hRipxDvHWgA7H9ofXZaPx2O3b5OH8zyWyQPKEHFold/ydAk
E530CDSn/mOqNo958hYJQ3o9XxoYmsTN1dha7g2COQZUgzq2VHHbqMqqBVFH0md6CW+GE/Mxi6w7
NqD0It/5h8E/U5NV71unIk8WBMdsQ1D56EcW3jFBvfY+b0htUfPuxwGgwb7D0u1UqqX6STMlDqYM
4BiOYU4hG0Tlwm7+wYRErllNPDowE6FC+MActkuUSKS7Hm65dAl+ptOgjdja5Qc2vds58e3CFDAm
4FiF+jv3dD6XZowGBS0VHqCvRdJUcz5o7Ff7OMrb9xakRd1dNmj4TrhlI5e2s5jjAZpz6yhmXkMf
8SkI7xPQ573KHqmfNMwmIqRn1unk43jdq5tpKpFlJN2S2FEWaoAgRhmutwfgWkO7MH5xn/TnZnn0
T8LlH9qCNYZ0dgw3hLncfxlSUOlqlZpVrsFrKqrJ1cj66o2igeHyQGvSmK4y7vDXxZT8C+5ZPOUS
IydcFEvTJEASh8zAZ7AZiVSS13y+cfmDv3W2f36ZKavxllXmsYQRhZFSHar115W2AwfiZWeixOYd
unrfa7CD3iNfWvp6jQ2omqcBVAfDaSk9JnNys9cax/N/ifQYdXdBObuL760iqZ86S2UcqUhbY98L
zGve0i7Q3CYeQ4Wg6N+DIUYbUQysAXY/xWIsj0mI8b5dH0kYQPYSfFeejTx+wm1G+wgDW7D+EFlK
UC4Yq+E5WuPjtb0KM2AX3jk7PNx3cx8HT+MPS3L82XIlDLKiCrZXczs6po7+smV9Bof8CnClN/p6
VLM/G8KCc/Vmh9RkPYzduPTl/csYL2/cfO7eblFdrsKVTkz5uaCht0c7F391fOT1hnAsNAvbVqLV
dv9ISyHA/3dOtre4mjy/lmMgh0OBFgyd2R7g9Kn0ybbcR8+fEIgrqwK6obUuFJzxopvDmLdjxq2G
IAcnWxVlD7fFgF9vtG9dWN2uej/jworXkSAk++3eoelPqkkz0kSxyZ2aXxBM+hNA8WLLRfeL1C9f
TcKcXbMRQVmC6HCkWwD5vLbl9dm03NjfCqeC24HT3yoyGRR7Y1WODIFb+8T2f3HXhpS1LhZ5ITWa
kRuyS/Tm+oqCak/OtNxxelvI5pG/nGY87fNwPG2IA+Knw9E37/SWacy6q+cch6WduFePjHAextlR
sOvKAfo42oMv8sipN3Oucu4bsjomTkTYMYX+X9MxDlx8GbX0S5CsMBejZ/U7UIahOTEOBsw4eIk8
7DTPy8ZvA+dosY1GT7zKGD0ddo/LpVAHitAkQRUV+WrbiBA5D8D8J7b16FC52vqbgY1fdaEDUvyI
lz7KgAowjquae7P1gD/WMO+9x2KK1I8aTgIZrJbcAzABWgQspOJ4I7TmLyl86lSHBmVZdWdIoS1A
BKVi5E+NadLjWt/9378qs8ybUPKEDAs0LO9Kyq22FyqH/149SlgkM5vVfK/1c6Ni3ENbJKU50R+u
HwnPRASj7ZW+EyjPO6n4y2qpYhcGk1zXuUxQekiO02lHJ65nkCDjlw9dx5GblmNUNc93FfyL+KD9
sDz5s8GQH/Jhk8JEwRvMNwIQpDHcs/Dl/USd1Un/8fEfSX3XOmGTQvSmBBpkm5HufruiddjiMipF
46kcLQQvrVZyeoFUL6yXI3CTXWYu0tmv57nQQfPcgbC4tHW3hfd8zhZTK7pHFqcW8q6NNIkOVjqz
wWKkxZGP5bAYLaDBpd77j9fE9+AG9huxIZrpYfncGfVbcry3QH0VTpHNVYixNuOgrF+M1u9tmoML
9t8uLDRdg2DeDLeWbG7zmOhuhl/ysPoeEOU52DwEUfwPHPEbOoQypcPbE9uuvjne4ykevhSqPTCx
9N6oOSl8px1kAz2ju4kiLhDUymA8+e+km/dpHnKX1hI15qtHTylniiQS9ixDwV1BpQ4XQDcYA0uf
YEvt922PxDKGe30C8uvSQM0kwj2CKjz9WXmuRZqf3YAHlCbjCCrhiur10gfN/TutzUb2DMjH17A4
kgZkDsFZjM2Qsg8fXhLIqdblJbkid4VrZy6Ml6SRqxbvZOMo8DocOUGyYIKOI8ypRAf1o1tLfH2K
Kn+euZ+Yd8jHGDUU22tmV+TjtDr7Wu3IAnFtgz1eSR6HMOer96PJqoyCZTYYUjY1FiA933YVdflE
6q5tLpOnla//pE/Cnrv+A3Y17rnxbdtn8c9lWaue0QNawN4peNhDRnMnA+7kP81IZmeKgHVFLxCc
ivWCz1lHYF5hwgJzhHtqh8XxvaSX3GMUFZD8JQCRi65XRZNAG6P9tDEcXoe6/58gMnxYJ1+Nf9Ou
Re5Lcqq8+b0pH27GorOh05JaKCJpCxX0ejlTud4e2VNLGiQfSJjiDnsBu2NzMqemM8hrrfCls3AP
u43bSwZVvlCZdlBigeM/RdN43Re+GlpAittAEzZe+cd81dgdcu0DB3T0nE1POFRWObtLN6UUZGxA
EmWFaB1r1/dfdCMzZnphxBsScD9u5MP7ed0ycYYWyu/TWsWZRUZhi3Zl+kNZHIpxqN9lpE99LvX0
fjHO5I/umMfkUbvRwoNgvsNpzJe6QBvPsIT6cunF5Gw4nqVdn2qdLXEvmFHn4vSPo/f1DdM1BDme
3JTO0B5Xo3bXR0loK5f1bf8whONsc1DZkcrnzfqnwUZGOYYxPKyCxKAm7MUdqUXlPqVxUwMPTTXn
/Mf957um79vqb4VqICOo8P8RHirF7uB76hS1pZTbu6mj791JnupNupiJswOhVk0wkTdS/fM+N/Wu
mGFHYn9efhGGFO9uNyorivmacvb5AB5439LaOfovbG1w3o2a4UUv5MGFDVQkAtPtC7UKHxiJfPEW
SzCtFZDcg0ztQWFtsQQB38LStHWrrnwYOiEmqm8+FqnAuDOowFeYKagcBAr0nxEF5FyUsZ4Yz+cb
UBwJPiOx1pODPe131IxycUmsg6gRK85+Vp+YLHzQN3ROPRe7SmLxPBArEeMkhEN8vdRUUdgFnQQH
WFoheyDXv3LvVTdI6lVONu/v4QmXDcsmhF4C46unxKBIprENe96RjRfxcPZ1gnDS+qz6iyJtS6kz
NqMB6Tl77b0W/tIHTJM4HovfXgLoyzpTPX+U2wTfffPKReEvIdGESB/6ICeV9AioVYTZE5gQYy/U
2q2PyHiDdshjXFwRBT0wNJqywjpKvRu0i2NXDm4MXw45EbDqnREKp8QYXwAs2mkvl/BjF+HBszHe
k1AgLtsLVGxwJh3yrfhq//PSbH1NVcdQ44HHdrqgqqgT/i4JkIfpkqtgirjXiejrzCdL0eLb0Zjc
d+dLEw30DaO+Et1Ogkl167RLbDt5T1tEI0RbYNdclP3Cvh1cjDNbDSO0TW4Ka3QuNUnZZFsxSP+T
h7pA5ZVtRAfP+sbmPPIBs+sV8gbTe0XQhdBZfrrFYYjiGvYX9qsJZp5cZyIhcFQ7HwR/u8UioBJH
AVw/gPAoqmZdTjBkrjsNmzMFHtsLJ3SlFaticuEH1t1lrPF3p9iLX/8UxDC81dNdUes7Dfb5vEM5
5yPO/AviSx/v+rx0VpIGkMw5qV5DXw6Vo90lR90jUjFQ64nvxgUmOWUZRQsyh67xB4cYlcT5Jr6D
5ZPPrHqItAeQm5CKxPbQaFGDuFfVUuNcxzmA0ocjLG6/TyDt+k/A667MlZRoYPl7GeZlrKV1+SpR
LLeR22HWubbrNcF1VI4ifJyJfTlYow+XRCuFZiFHXmhuljOooJn3Jd7z0Kypu89F3VCJT5zC+yK5
1Vo2txk3g13lgmUoUO4qWtw6+KWYTLWXx74tnmRCDg1YLAEIcpGh8Gsz/PIxYt9SngRtxuOoiI0y
46td3+d8XI4zkSbuVfGoVnCek1+XZOV+sS1JXEgko0JrbB7rFLOiw9wfnYKIywOQYChmEcNZZ0E6
8Kgb4zPmjrhzrb6OfV8GjBIZ7EEwKHt9atkBur3Tu2QPNY63OjouxqAStPThX9OaPGgWRgOlccWu
Gxj3Da2RQiRR8saWaNPsrAzHUaaryO2OSP3KoMGYw3D8MEZhl7FqTN7tTXrJxIsUnJmhDE5dGfYO
GD18nZ8RDQlwNix4m4zR0ipio2ik+UpoG0bVF2RZT0xEckdE3sCMRb8xR42TMVA3erP8V5dwD0HW
cz66lrrhD+ette0fQ3hMGolAiDzMvbJkEZIJHPCSVM8wJRSzL+fGLDyiWUxxeXo5/vGvSo17bk8V
K8gVx93dzAp2dBYq2XqjINzVW9l1seSniGSWF0P3Pq80f5q/TfY2naPO46lwkxpek4nzkm16xlfs
HI3XfovRWeWZXUGFH4EOiFRKgF6WKVGzsWsXlzvqYW6LDEYBipnRqiG9tlHQlmAOUWNI3d63H0t2
MttMaRiMurmbSTjlub5fsO00CY9TpqrnoOtGVsDZeYiiLe9RzyE71XW9DYRpjNuTRUzPZmaB4kbm
DP7vermZiqtpz9IWxJwpz+ip2pp0FQlEKw7Ub7+thBvUu2bhI9O1cc+vPNmYXvTn7bWxB97zN7p/
qYg/0UHgPR7JC5y9tkqbRCbSfbtJpDySxn0NibN7jvxeDsMw40+4/jNd7gNpbgVF0Q1sHDq/MQ50
MiZfcddstWY6+j8xzVgWCH94H21b08Cl8kopuvrQfg96mel0vdjGdSo3+hBiKlab6rbilb5VawoA
SFovVwO6+Sd0CJELsF3A6hRQq6ABYQnSQfV3Fcp+wrIOP2/2t9Ji5ORD4g61/HSA5yEIMUDeXWtr
m9rDObRzCpzVwgx5GM90X+3MnfqPZfo+3m2o700rJytuNFa4epnXPuKr/Ic9bW7uFamq98KitIWL
gQgQVpCb2KpdLxLjjslhpqfQdU4ylBPDSNp+2EX7pGhuE3l0xw/mS1dPHXGOQnymvi8T4g82qA+e
RlsvLBEBPt79cbSrkSNolPHpgmf6FFiXBcrnNx4CiiYLB1FsS1kE6q93eUS8vfGpoGP5sijVMVYz
3JecjW0CG2tyguJxsOq+1mEFX22rHl6j+wqwCh53Vmhndg41PQSzzIql/dJ6KoTQzkhsUli5doVp
neaTzmk8hT5MrMG25YRQs9YgTMqkk2MvWjCaj//RSs6cRBbLjiX8DuFQR0hnFeT16bNZHoem2hJV
jyfvGRWeidebY9pjPY9FYDWs6Fu+ZzeW6KeGEQCAxj2GBLDyfaxAAtIwItp1A76w0w7ElKIG5JMB
ZTxvYQkm15hoTtI0WKC3JOKbrG3nQdDR7/FW3WZju16xOE3mwryDxyrFLYsb5rogZ8Nr3k1R7V7J
snMhRGgwLOG+a+GOH9WcLO/kga5MEEaLHMb+a7i8vm/7laBkBpOxKMn9isU1HsBy3W8zp1fV87Hd
mH32gHtJ7vPnzMOR4INvGlpIZrv2284BAwwAneRof2s+zl/IGPlhkxnnWkIcDKlXuXYLUZ3MxOEi
WEON9NNGmAsFiGGyaSVAkpDqwCtubToIIQudqT4CAjhiToKVUOsDlogl0Yn7PzormPtLTLqxUIkK
WDniMoEez4HMNYtH4fdt5gN7YyDuQ+xfwbZYtEsl9IAw0fmoDPTm3ahu2L2C+ft9wlPh5jXl+b0h
ReytqyBqIa9z7C9T8w59hYf9nG0LXvalFGEZNmx6tRsmTrHMZQ+jrk8k+1DWtARwM5NPeZAGt/2S
l5lsNtgYAAJXSOOj2+zvr+X7myVQtNn2bOGkTpUOAyTYTv5gsgXh+uQxkzR9Q5VZqozHdkVhxXKk
tRYBwLXxTefRDqp9U108ow9oN0+H3XF0PxAJUEJ30N9yIh1uO4mr8NQLRKn8iQC8JWe3M4eWzg2v
/z9i6HLK34ZualAQ8rDH5svgi+m9hD5Jwf1oDlfoqxPC6izW6xuRy33cIsAUXsLWTOkgdpt8p1Q8
uzdiWwnNSENIXcHZhmLw3c/QDkCK9OAJP+jggeibu3euFx7p+G7qQt5c0PgkFFKiuJvUnXzved5e
Vj4SoauLeMWPQCloccjtgap123dA2W3iEp+Jy+vois0PG6UlYCbtbCmFUMMPapchs3HUMla+9O3L
kn6uBqfy8/ouAodVIFA+cWUCIwkVt8ylo0T49MMR5Uct94bZd71JmJDGvUf47/yBBzxrKZ0qDmXf
iZOO40TIfDb+p+9DMQzgjTgaz6alJgJJrFjlaTayddDS11DWltlKl9sd4vAB0QPboi1eaY/t/g/S
qE/NWZdWTrnXrAMIuWGiofaSYRxwp+N0Q1YYNAwFjqMt7VqHGhBfwOrB9TSO5Ats4zUW3xGKHIE+
CYFqU8MsSZtXOrxZg8oXffMYgSOGyzCbWkN7xR0sNeVpqNwQLKKlZizNuhd5B8ZAR3mwU8Y9Z/Zr
vqSG0DwWFP44UV0pehLFtTyq4TfeuxXdev9vK/y6h0vIFcjXN0jekjvSLIwGTIrZW33oLda+CK0U
GZsLskIjmw+GvDjyybfnl74/+rLbA+d1T5ctynCPzhISo3Lbv6SUzmtCI6ny4yz8jhPfcxCFP4xJ
fi7KY8bjEm/s3w3UKrvshUZ1HcE/AQMUZmEs4hXqUJvgpfy4X3+2sgBGwBIpPPx39f1hlO12XFU6
DRYkDP2ytq7pLY1hl/Mblw/EWI5zPFMgbOy03BGKvKHX8NwZ3ljFmUmHyGVWs9hjNWKzRomMg+Ji
ybm/QmKlsNtDcM54Dt8eKa/sl71SySTKQlWRTCxr9WAzF3nuAn0oSLWfaOlXF8LLkR7ACXDKNJLo
zn+Wv9HV+fw64zYwb8CJguxUy2eZs8yIYLst7cx7we7bh9GsSQvc2HLMCMKqayYbIoa0PMEdsdkd
VrTejPNL8GK7t6IUHEe9knkNntZTd3QSzR+o97zi6CK1RgaPMTtlNXvxMeGPGXTBQ4gBSX3mX+Kh
mUJ0/eb4Ga1Y2+szJT/3kZupfD0g6uj9FICDEmYb+FHjw7Pxtv+WfzDZGvdFLDr0g97dCl3sCGos
R1adiCifZyHmPM90CNcBYyLG8a48D0t5wWBEjxB/21oWffDTZxsOo4CYwZAHVRlxWya9dnr2zDCe
J6NS0zdNfoFE2ah6EgHMyCI8m41gfV+/MxXPe3P08HaMfBW/lR/8mj3nLUDj90sCVymRVfKRGGsO
+/MgEbZjygQhUzPHQZLFVlt6Q0XY4kv9fq89hXt2/yPCee/rwisYn2FFrvECHTSfEt5NagZX29q/
ovsEh2NFfdFGewfQsr6FZRVDTjgx4/96U+VOc+xMo8V7yKpCuNq0W8M9fAd0wYsKptzZpYC27jKM
1CRuLOlyV5XEcnIVnDK4bkXbl7Dl9m1Bu0N/SfoFj5JzDPWX06wF31O3pGJefJNa3UZbROsdIqTL
JrvxBsMEj+Ar6JRLkCKPcRZfJ28f3++dwdGhHubE/hoy94I1sXVTQ153vF6EIfHmUUt0BI2rY7N+
4fgDfyE4eEQaGVtF6x0lJ6MVSm3UvoGZHZ9uz2WVZ2nj/yaKHfYACFG9bD6waA6j4fGRJMDHLKNW
nYATJSPG84tMQdOzrtpF659+2K2qm5LR3fCFxJdKlFn/sInZ2Vq9864HgUvePaOKk+EUegKH/nho
gZKReCN+fvejeFx1D2R434WJiA3TJFGSUtSI7VILJ4GmDb6Jk/QSkuXJp8LOvQv5DOfVNQgo5xQ7
IPC2cMN++aXRPLLVG2FyHp2LEC770TG814cM3HcmhK33ihoXokhAKyP8jgxrrYXVRt1z6KMSPahe
u3s9zN0ugn9MO5RkYysOdYX1es5LXF4uVgcCr4+g/CbOp2ADH1RtqFIYE+uT/qFg1WMgsFT3Sbqh
AMieFvUPfBaFWKtgrh763uVGsRTGlSyoX8oVILi+AxgfNinPpHhBlfrgz6zkPlXd9ik0cUc51A4v
Bdz00NNPPWoVgyPneOVtYMKRnL1FeVa76UoP9q/SH9kZmobPD2PE+xv4EaR6YNvxrtbmubspQ3cq
ImwrReGYJPpGb6BxnME5p9b/OwaCp8CzJngSBjyg9w8xfkE31sX6wYTX3cGOhc3nP92m5RBSxpqr
UxX9WPHq3TrCNyACDjGbWfjhmsUJ7sGFbM7638GPPgUTmp8jG7FkyfbUeXry0aSLPPTGvIFZBwUm
slX0X9Dt+8hzrcAv0hqMfAovzvxIosPPO6FWxqXAk90Fay5gFCHWY4xDRFzZRDfqtAgeqL2FXquL
W+RE50AXJq63iwoGs+FfcsRqwDXbHpXh1tu4CL2o3snqAxQapDMk0PvTrLgVxKEY587+ZBtPodlw
K5nJ8liybhYmKm3lAkup0k5iTywJBJeQUsa/U+8eZl2fnCleEm0dX9vLmo0RB7xlsficL6vjKrVy
6r5WCELy0VKS2o7xBn5sw+Vp2q6xItANfz5MmXoVZjllGm0sNPF957wn1EXts/SJA1yGmyityp8U
HosBaShVx7PwCRBH91qNw1e8zqEh7CYtq9+m8n+3SdmTbbBHD3luRUEVetszohh5mBIumiUu4xdD
m16iTT1rPZLgFTipzRRnfjGjYjuDJEkJPRZZC/SrON84Bi4L+6Lurc5/HhOJi09kivicMsEBjuYd
cMnsFa82t4uLYdqypuQ9m48EYjwDg9+9ejuH4ZfisHtBr1axJcaJQdEeGRjJdNY2l1tILLcI8bhd
K1U56/l7U9qNJPIYpbXc+/CoUR2/4Ea6FffQMirDeJERP9Ei7MiWuVsooKZ3zoTaAo4mR0XP/c+l
psJD9JESABVw3tSVTguTuHLu6veVSkDV1f8reExfUK1luXRkPl5dus1bzTkdUfqcmNWuJIZ4+TjN
YJG9kd4B/8yl7ymwQ0O6R72N+rMTkmXfJ0MRNfQSAPT/sqjCwLlpgGOefgRk/LV9ZUiZejI8OqcQ
K2Wh98c4jKLKDlYsluJRirgPkxK7i8kiMjL2Ox+DFuxu7xCFl2FWPo63QcfY88Ik/FhcrH9XY7Mk
5Yqq0i4Gq8A63gcicagny63TxDk4T2t9SkFS+sEzWdMmqEu7NdSCqRbOzA+jrJM3/JXh0Yun+KUv
klWmpr6zOmjFTRJ2y3nBQxCy6fhSGnMSNAOjS7UO3OKWys/SDmefHCsDjXfBiqydyWmaF8ZiBaDK
fwm2/Fq2p+2U7csF1KRqNFVE34YL7nT0jAHF1zLp5s9dcXmQeM6kfZOczX7CMgz+c40KZFc0dHto
yo9+ndTC9VRST9bhvb11yAOqGe25jZIJG1yLHJw3EjLGwl6jHQCioLu6d71K77esdAQi/B50iE//
B1Zg3/cHrv9zdM2ciDF18IuFyMjB3e37e4FE+WKqYoDQbZaTK9i8krcg60OthJ0IE0ScazRf1aN8
3VJRp3WUbq0s+qg8ZaEfhEs5zXk9FuPIO6MBEX1YHPP1COdbXfBhWE/9/t8wSzNvQG/WKMCC3c8l
4HMtFrGPWWUtaDMVLWLq/x9lxTfBSqlSA3p5dKUFFWw8tEQuMLeG/GpQwREM5onxfn0LbFjs+76j
cfZ7hm+fnrsAX8kp0c5YAqEhB9057I4h6bO6/6w62iRQ8DdsfxvmbqVV6DzgCV6Whe7/cLPXNfBG
jfAoNWdVTyA6I+GhAq6Rds+DbjXY7YamIlcZAEHLR3v55xRsSsa4HoLLFIn6Wv2nF1SifW7FmjAp
fM6Z2HqoRqRyjvguvGdz39gCyTitTObEUYZ7lTtB5gkxVM24Mj2mJsNcjtiS4St8SJKocVn1cqIT
faWEh5hzBhE5GN7Dh4z/tvMO6B5SMg5v/gkjCcjMFozd8srdsnsfKxOwi5p6jL+V3sXYMZlG5OTL
o81PQfMVGNlcXpfuIGY19mj6sDvphSEFUcfSp5L/FQncK4ApmvXyNUQF9hTUCDXSmDfq38mwrJvo
zetNnrZoSWaqe7YuWIpBaaVvBylv6LD5CiPBNMKswXpEvZJfj+gyc5l+SMWaWz6153HQk26EKdyg
N+Ekt5utWuSCHnvXDML0/wF/7xO8yS90HTMIjbiVzy6zFsmz/sVISI8ZDKED9etNZVwPr9jTOuBD
GDGBdy8anYOlMK66NxZmbfr3P8tu1BaBFCjiJS8/vCu1ZSG6opjpva5oV99+ZYPuWVV1wDww/Bxw
JhxLvMvDuPHvlmj7Q9se8HEGAnrzxMXrJ4EXx6Ar7h4lAaAxE7Ascy1JSn2EZi5j3QAhuOXHnnIx
m0jq09RBoLhRk+JOivSxFJD+3534goEZfl8Mym19l+3z6OLAb2pcbX+cqg6G1GO4EpVZ8/kq+Zzb
Lk/9LN9EWJ8JxD+BTHejLQ1J9feGP53z8cUbaoWZwy105/Cetr8yEDkSUe5aEXlKLoXVqRpJtCPI
Q0TSeFqoCjjgqa6mjv087/2X44YXsebD+Qn4AwI6iQtlSedWiy6qGjMu5NSxEIXyW3T0gVOZmoYy
9ZiDmfoVSPK9s6l00NhDALQ9hhBmicvSUHAYeAV9PThRwUh8G0HGpSCKy5peppMhgM1scFMuWGeq
3A8EK1uVPHFqVdUTV+kj3F4NPe9h2xcTwTdOklqkB+PiKN1kauvXHauM+1JgWFwiRkSsLbTt5h/T
USyUZ2xeCI+Lmkc6eemwCmDLdgLkTqlh8Lf1j3W4ys4GVIaoD/0mHxNFbAq0o1RfRKh7K+qdveEV
IaBa75HEv0LBgO/HK1fZUd0IjVQixu1VLj3Xu68oFPsZnrPKV9068vFdo+VJjJQC60TBhli68yEp
JlJ9qQfnGPpxfMIC2blzUrhtQRxsysOy8w49PURoizwqA/3psRQFmCRzPmH1Gk8ecOsrogNPiNDW
UMq074dfWG6wTLzlFUg0qsz28U0wNhsvLGcYHqPvmhHKfVG+KD7ykJr4mzilqS9S1T4t9UB2yfgF
ZamWATXu72yb3Eiqx1cqVwLe/+QWbtwokh1MNY+jef2alou1wYg+ZOqzg9W5hQwpscUuFhMHoeO9
/LBwAda6eqQQ6sThqJhpSbeLFIwfpr45qRgNUoL9GPVw4/FrE/Z+HpoHoyttZaC4yhfRFC51zn2D
mv+kfDEdmAk13vbXWXQsxJR2DBnAEQjiySk3+hG/PlW9nWcZ4Kk2+k5S6JBdpSYNRVVEbiE2zC5w
oJp1M7PdE28BoMry568gGjfY6w9QG/9I7n+cGJcsv6n6Y+RA3i4Iz15s3pRgqSfzF1VziIryps8t
U6uIH2cO8fxN0W2C559VZcSbVHPxC/4sZU1Ek6aFv9FE9l/E1zPLhl17sKRejslQiMGEUp+d9pwA
e0iXsvrWIjzA8/0tEKqRlMT3UYEJtwAOjhgYbR5dzeiSC2eM1ROCq61BpnCFIsUUUiKxziXIrnNM
K8Wr2JYdM9gmoyHjDq10+N8f/BHFQ3G1ayT+cXpArNYJKMEnqVH3LHPksb9qzvps9O90V5MWL6cP
khbEGQX+kTs9BbT2MLOev7WBMslj7BH02OVAxJil1xWi8LhTmy7kVN7XsbHPkonqcOH6QbwMxz6t
DfHyzSAxZ/7vzENWwMb8PpNjzHnGpE1b4rzqQctzyuKcp/wNG6jQsJJUjmlPMPPYF9+5kealoTzh
bKV3r8VkqlqWW4JjGF134G/9AVppgATrmCiU0KLpnSVIiMp7boAPOh4xWDBbc12/mrylD/Mn5mHg
FECW13scK7yfNn/frcEXGfRSIA2OFssyE0l9sC3FTUCcErXLo44XCxLeyWVg3ztn+66fmZDWOffB
1JohyknpJU4/JWFEG6MISzm8IlN2tVjiQAyjtLUxWaCxBcgDYOo1W6g+PEWYv+kkI7c5pnR/7iU3
nGK/BDtIcOpje8SG/Kn118FLV6mHIZPmvK9Z+0IEAzkRnLCC7Bez3puG/0W6q55fnFvo5x3jXuDx
ztNwvx7575GtWRhwOBYEc5pIuaSgiTvH//TXjeJve5WuuFQUbokDHRnQHvUklB3LDclNbak8l0Qk
1m0hWbMpWTz1AJMRU6koqZ09YX5TiL0zmNVO4hRWwUGXpxxNc/NHbloUuQsm6eawma8R0SQ8VgOS
Z7DUIIjdxrxpJvzL49o4qB4IFmZl1N0/cUnqCLPIn7xsRTRZ6LJ1X+6Gxg98uqOQQ0uet3QRlKcH
bUVKbNRggRVifX9gMk6hd90hP3stBeuAmFbNh6AiuIKVENXs69leJKYls8YdFc4O819C6tDdJDqR
0zVSzMpeAXQd+EIOChv+yvWUmoXYjDagQrQ2j1TSMGLMNbY+VZ5R6nzYUV9+h2/S48+EDIbkAFV3
FtKcQ47Ox3NFKm6tLGxdZGXhSsbX6iI0m108OEjtvFSE5Xl8CVQ4q1tEK1Dpv8oRS8BAI4n7PEep
xPsd2rDfk6zWe8t6k8fB4v0i3GvsSS6WdJK1+qDlBzAWe8ylZGwgcd/JnreCNY7yTbBBCjqpdodO
9WhhAnAtU2YRvTq2+pmlN6BveuHvNZzVupeWercZTk1+CFLWQ8KnKa+bdilpkUB0XDnZQRe7wzfz
Knfhrz6A9aSLF09CncAuBSMb8wRTT2pvhlsHQJs2vaYcePJse9Wk0OMLui/R0yDEHf3DyXnkHvZD
Sotti6xTpqW6ofIuMSvjZFWxFpEf/sH4uEz/fXvqboW5q3mf/hVaKBoEaqmjeQ5/wTl5gNF0lQDn
hGj4v6/fcKxCZej71WND8WEI1WzeUcBj+qU9+RKVuh+iRpeN/oa4QAOX8FE/JCjj/JD3NQDCaDRq
TAP+krBwNeWP0zL9VqVuQwH5Bl5abfRy4hyMdzlnLwxzjNkIwnu0yJ6BPp9cpo0E+S2VKqpRVpAy
g2zbruTWI5xWaBZLKI1rlykd49JTh7bjru/RhCMzNObT1FUCnOWoAmtYteHKeFs3egVnDwVhxUCz
782BIDuY1Gn/NAY6NKhLWg7NImcJ7Mfz5eL6KfVuqtZcazm0aAgbLLFs6EhYupL3jroHyhW1m9a5
+tmqDRzTExZeplsSqbS4RLBBuEKSt6ujCXUcKOC78slFjP7UIKziexGvCtyVNIulhFepnhlfKlMg
r+1VR0reFJtmHsVBb6mxd8utmuKuCU6vlXs9Ec7M0ydyjmndl/eK6Rmz/0UqDdvdHTmzxyl8B928
5cwnyaMm0ZB7mQewnZD99/QCxfIqPDfmammDQVBrlOuEHfBmWoyqopG+en9nEQpRGckhsS7fg1G9
lcXfpkKfOzCaL+I8+jf4+KpYw4efcpZfK97xlM4Chwx5AGxip8Y+RMR5DQPfkEM/xsmM4qpIaBIw
mTEgyiU1E3+iU3J8C880viW+XfPDCN5i2649oCYz+zejvtXmt5+yihw3f4tl/4ZpK8TDWpHnsZGg
A6H4jhQYI3zVFU14V6vhZruT9I/RTZGEEgpX3aKoqupwNL1hZkd+pIqL8Z2N2H9QafVpkKjeNtrX
/2tRKctWy2wzm4d7A+twsRhQdFbl7SL4RkoR6mo6s2U9uaKg+Bnd71gIDHpMqJL0+aqk4UDz/KTK
f5TZdg1WtsJBjWdbH2j6NJJbxzNiQC0ixqXuBf4hBb2dXK/IVG8PZNa4wvvMqdyWK7ZPhhsva4wT
jAMRRr3pGDUt7fD7LAU7+ZJeO8zjSO5ZpkoEGrE+7MimCNzRJLH2HalwKAjAup3uO5rOeXKUmTWc
QMTwFK7VgPmGYaLhL+qukFp/SJrN0+Wnb30q8WFe6jZYbg7zWSUQ6UbYGi+gOBO4O4ogusaUHQ25
k0NA6T8GUjlAt+b6oas1tZnOiLwvJQIKrtITZBE+OOTn0PPqLk8wQlRyN6hOlsMwkWlvsCjZpPb2
Ex5eyNhAM4yMehSjjwnYlwayPA60uj4KlvdqBfBtcQA6PFFGyrRgeDtmmv817Avp4savu6RHHSWR
qpnGwMBZ7hDr289ATj+V5uQrdwjOsk41Zd6QGu/OybfDBPJ/xNWHnkqhhVneBrHQ5K86io/pfv+o
qHLQYv6KbcvINvRyyOUwOQJDtj5X6dbDV90bl+49HNic+fGi9uJef6+tl6pubIMsVA8SEk9kDwVn
HauwBGsHsLBSh26nz3CcJkpLCCVPSFXHJdABGvxjZOAwBU61ApWMPXjNNUPjaBYc88B7XzjgQnU2
QiGYmP3saPZiyLJSPCUumDY5u5GmHW2XNQjtrPQEui2P5Zloq71ZJQnaDm8XiPNRhy1eS4+9Pk5B
odIaMms3YhWurWsALGl3jE7ejKh5o2vluqL/L9mg9lge7NdMNEFyb6YbSFFMLoMDF5Qk5o4EmVTO
lax3fZSJJnP7iJoi9XPEiyemOojo8MXBXTGTtKP2okEa5yI2s8S0L2DvPjYvqFVxbLVUqT2ufN3U
riz3Gr4cx/tzeVnCH9Zedo0HmffdQxcNLZ0XasqSYuDtS1h4WEP/FEmkorTQJPTXkkwOIrsT+rTo
br5QnaYcU9csZdpgxoXJN7/5UzV4B6yCm4DNk3YJkzpTCy0L/Sr09e3UfQOAicTFTOZZDOLpH/b5
NhEE9qHGuPSifg9hOSX/MS9jcnKK+frDPXYpHCD96kFwdsXLwFXU7XFxod3h5wp5pPK1kig9Rpox
5+Jrl4CEIzbByAWf/JDNfooaDRMl+hOqRWz2sZjf0Xf0oJBuFivToA7X4QwU5vxVJV007tzE/8Ny
1I5nzBxc9JOjhFI9KOF3CX5xswvt+kiC5lKpEf17aNmGO5n2Aj0m/c6rSuqu5Eo8x35R94x0uzFN
xi2M0Qp7bNCyooMqwREVXJhyO5jmpWcx7pCX+9xbaiqFiB3EX9kZfguhD4zbw2nHZqdN8Yu585Vp
xmdGkwFvIyzAMXmQwCksXsrFk4clLZSSbOPy8504Jrxyc/foRK3+JMGSEXznSidB72oS6bnAL0OH
gcNLr1g2P5AtLPuXmPaxv4t81E5tKmGXhyRLz4P1JMPCfYDdW4guCKwL5ljusbD9VWqkvSCQ16Nz
3vSPU5I3or+7G8PxeatE+p5xEcc+339vCxjPuBYvJnizOEU4LU4hmEIagXfzPrJsLWwFsiFaJt2i
+FPkfuXdfyIE4XWDVGUBpq6TaQFZvngTGM82lDiKvvlO+P/7lKaULAIF7Dksg1w9f1fn0+jjT6HJ
beSjYlYxXSIE8CLUyS2gbZPTanXqNPMV0RSiqJ9VvDROxhPeqdesSIT4bqrJRy8gPOcrXb6/N/pp
Xub3PHYKHNtafzv54fdAgIOUOKt5uU57+LBH4t3L4kaizEB7wcbCPv6dHxyclt+SUYvLf6otXRXs
SIgDvVbeA9YVb34osZJpSuHIPzFXn21pEzcuSxvEbBxg2bhBG4y8mm4a/bo4S/92Yo7pmmE8OduE
Fk5+2rDQ+TtF7twvcQYUENceyUlyN9bdbNPcWJyYjTdUXyD1EkRQt2GTOSLcST0It6XnrvpzexSQ
YRlNbgfYq2siq2Sp2nnsjE7hiewMpZjk8TvKsHtBJ1l/xnpb/l5jdZN10le/aqDtNxrUPPGx901S
iS4P9RMxwT6VXYIRRpNfkbWoRTyyvtGpzif7TB/dMFtTbpuZenn74NK5haSkP0NwL55JNJ/tdOW8
0eS6NRjQgQGcEU53Xm3dxepqtEtEGkTYsuZpNkiHX+rdkROVLlvQYPCewvn7EDJ29AHPE4WHcIYR
qMMu5yWVl+3baVTXm3fftdJa97+BWf1tm4MgR2OfgIlpA5z3LYvg9pzU979qRuEsYdrDuD28Dee3
sA2nheJqBc0oTF9HJw7P1W6+h1T9zIU9heUGSHk82vxxVR+7SBxId/iZA7ho/NkaafKCkpTOHXuc
liaC7OOOEYTsNQ5jja7MyS2/8reGAKE1LqqaUB7NB97tcnEKHTLkwbbynDY5Bq38U9ZnI3nZOWOo
CM0ttW5pcJDs8YfjBFYaUWIplm0rS+Ty6rfq6QetrPqjeQvRdPSWvLRLQOzOSE0Igc6iA1idxwdM
K5P+V4qRFrWPhFFibO3cRaKUt/mUXUG73g4iN+GcGQJ8h4Kj5aXj5zeTNBRMp6Ix8odypW/NdImG
6/iHX3Ik/g3mlSXpJrhSVrJ5wbMMftBu9w7CB8uOqh0YDudnrhi3oZB+xvStT/jK/FGELJhoMhYi
of1rw6PKuS3HYki5qwD6BL7pWdhvAm7qYVCy1GSPPieRnUcs39R61E3/axvSGCpIOxMVMJB7T9Fl
VT6YRcntwl8N0G5aHaY5jUoXAKSCFo5JmTkKaT6yfsXbQmyI8dwwzxfZYtLZcpL3jnNcoemzmal8
HyQUS+n62buxkv2bCiI77MTschk+0UPFcxh/r9w2PP4iDVOJdylgwIL9HFmlMZuMjceZP4hAcxnw
cVPLDagipZoP+tRkhdwYXc5kSPO7YUAg2odlzyYLlhM9S3u8IeKFBaspLY3CODLQ6nXKH3QcNcLn
/xKb+mfEFNcnxm6uC69vFkdtAD5l8O7Zbp0Hvpkq7jpN6C2ZKKSE3KTWOfqsw4tYFDQ0ngR6fnAe
H9TjEj7dwyW5QGKWeJf1ugs1KlNkzrntkg2m5p0YBAUjMklx92mckdOapyYhhNTOqA1aQkx7rXjr
kVk5M3+PYta3TQIpejmeh+GIKfcQf20DGdJM5VcUMmyn/Nh2+dD75giqCvLrUcGCH1EXFM1j15oS
PacDHZQxvTS8uZOUCHvpPvs4H6+2OsC/mDCnS7IXW3m5ZyP0c63mFUaohIfW1iaJvZZEiV5BqGml
YWg3gwlfJjfJ+OYoUoPsHnGqu6Tn/gS+o/ndTx5skq4SjZcnK3Fp66meS2iZxab8kysv/Qj3J+WS
iNeNN33wUPcr5mTa8HX7gOryIyc9IT9WiE3xIU5ooQ9ZOto9jR1nbk3jGG5UMqcZS74tjeQTlbbb
Q+yiDE/O8iz9YbREN2tlUXxaIJ3wYVVvaoB0TsxHvYX9SUePI3Qe8ccrVeLsr6vDCpDQtylk4xry
nG0vYsBpQw/Bz8srHKC+SV60Jiysiptj7EQBFfkBvzfy1sxgd/CNjxjROPV8VOdyu8aP78mSqses
W8CYyZnC0fucCyqKldJgfm82ZZYZfODhGTuH4r/mh+WXpU+Tj6/DZVfPFXZBkG0ooKh1wireRcBO
gUyAiyhqxbGP/Rzur6yYdB9rQw6nNqdvBCcJ0iDLX9pXKEeMIYLO8OFGPZ3AXN+O1aav6Jl8fNpz
JyXE/9lxF2FTdcnmQL8ZE4lgqgZcBK8nWnEP4tpeupiZZWGcohwj2V9XTJKB8J9HZGmxzwTcVgJa
/Rbi8sAPkYIMY3PBC20MvWU4nSEkvUd3I+CUJk6KoRMTlq2tgrgsZv5pywDlAyZSO/T6uIXbMYGt
TSmEB90VagmlVN1rDiFFugs26KBl0eyTceMkHC/mXt6+NgeGqivLL6muKATwESbRZrkgGLo7i8/f
LA1CjuBQpGNJrvHN6TkrqkjOQnRkEPaiqaKwPEEZL47QpDZIsh1JYv+1WpKU3tNOqa0993SX9U6k
CyKuMgFsnGrCBeypyAZWeNuIFah6kdpRGl1LgiNRGuMgikDQNEay0XlG1omHCJggK9yaNMMe60Qz
MndyokJxKhZ5PdtSiV2fruQiD1U96be5nkBEZNNsJyJcGe1pZJUy0ZdAENZXDexpeDbHGDj7s5ZM
/gnOXAbx20WA7fbqnxAk8StHn3HxGUyisXZPlzu/bh3uSDH+4xqDMa+5Nzqn1gEDkQOwWYci3wAu
sHSraU3ApiOmAIjmVE4tYtweDH4IAGpC0v8P55/FNOyB+wgHC5zE0I/jKDZEMpbEutt4fXpk405B
CkOA5egnRFTy2Kg8Xh2z/zlHB5V5beD+CO06g01gvfVXurCtVMUqV2c18LggAJn0Ix9sYbg0bkle
AS3JALm3EQFyd9N8G2JXoXscYDC4rrtoQWO8QMo9ZOUCP7SUzqPFVVZYPXQD4uEoB/AXCnRzr7Tt
R71G6qoxM3L7n/4nZMNQSbFgll/+yCYpMpb+5wTwZfiI7eoYHctIcSUAM+/XY/eN8nr9yIU6RasG
G4NeWy3bL956coJKaMvE3uj8nVPswfqfcbfcL9AJQGjYj6luInBZpjxLT+/lOQNFfkoCtpRerkIf
8Q37YbsUOiBPSsS+XwIK5KFHWZ+WSZ4eIf9NVG46LdtvIUIyxKSdb/uhhMWCzzMpSuiQHq4hN4CP
8Izhh2j5gVHFVnJ3FnivbDVA1Cd4eeLJB83DwgBVJ+Ljd3ufzjQoJyFh3JCAismS5Aj680eM1rHL
knKk/JTa/2/acJ6pm/U3zBwGJ92Blx54unG5DDDGKaz+PKJk+rXRLTBo8i42QMXC1cWj0KLWEdxY
joirwNJFZ5GMnWtD/26zCQAdYL9PNmDWgZ7bNbxK+KZ/kvUDZ0/3VtkZBdfnVv+xQPK23hcCO6J2
B2fFUBp52TAn43tuODx0Hg9DKd8AehV+Xe0K3OBamnyo7OvANW4V8KlhgX/lE9tVA/MmonGMVoLF
KgG03dHCjBuAzqS1MtnqpuaebknumCNd8k4V3X5xrbGqz6lvIwUkjeQoIVA19n1X2XBsLuebmDE4
sPKukW9dmubnm4FRIWKIwsp8rG8BeJx9hSCl+ikUrO9TGpHUnMQtxeFpGCaGv8MUrZpE2VohviZt
5UgFHyioqRsdkLZKFeBtE5grd3Ub3CGlav+uK1pacFFNIJrxn8VZ4Tv0HrT45DkkiFS5NShnLWMf
mX7sm4+Y03R1AGRnsWE2I3SWE0+96mULxL/5BvxjVi0d8sJE6qU9nikfat4NNGUDDQM4vsmwh3sX
r+XfnzfYRnBFC+tNUHSqYCYWAhCbwFbWXa6Dl6BWsqYhyeVPXT29UspH6SIFMDADjgXsnHlR5YyU
M2yHBHR/Lht6KpWavcNLb8BYSc6EKs8VgthIP0mMHhClgm9FGqhy2gY2u+9X1IXgp0KJTnMmymSo
AY/MbzZahOm26T8UMjBlMOE2KNbAbr1AOXB56Wdrtfk/dyxmCgWmgqR5Jv6xcX+MVEyfgtM0g9Fo
MVJ1On702XLEfwG2mLowW3JWYULWcSmo68eKpJUzdk5T6fzJnsFwMNFP5ErZ4T/14I5COy8rgFYq
MDqUYjvjjL18laB5/9Xd5o4ldeQBoQ2Zd/To/0z9w7Ub72pP+3EHsr4wWCeDV37tm9x4zUWTKdEa
AT0Mgyu8dsQqAalaj3MsIdlTsRiX8ouV9fipgJuAGXonUHQyicq/fhezW+j7LqDd7PxEdMOmcFBV
bxxn+t0uj1hfOV1JnXhVRxwmn0a/Oo5khygfljrIwLXNMbaGO18dADFLvXfGBJ9FIEjh+92BivIt
HbakIFy7qZyRTclkgFXIsYHhznRjnAbzqm+Mi9+EtU/i3g43v++/6de/e01sPORX/lAKNrAS8YB8
ULOqlQj1cqnwRsUlVaGWuXyNuDkvmw7+pD5VPryBtMmaObyf/IupkvciT7magne2I4fPp6cPgjMX
nbr/gwJx9vmk5eG9U1oh8w1FVQOtep3R0NvrgvyFAsFm/nXF02CXk2d7E4K8lwb/A3Yv0JelSUCY
RjTNikX+S5Yn3/oYs79ELlkYmyr2Kq086gUOxikw8qfUdcLQWtH7X9EpR4PthASPkM6rCe2TF/DQ
cstEsY4SLyVZ0wu/SaZp29pAnXS6Aw7nQa1/Wef3BM0gS0cZD+KyKZg2cMBf9SIMYxjNYVeTesmU
G514AcC3pJC2UUOnSIMkVIGi8K+G5ga8j2pHmtfXlXqZH2e1Mzs+wFqSZCCV/WVYIVQs2XIRhCVC
ar0ElMz4NwpXfQEjZRVzQk+W0te1KybKk59MxuNaRh/XbR6necYEiV2AYxogc3eE+zetFR+AIvS/
RnB2s3836c1ITehjN4a3Ur6siwBzDrNSVmbjrt6waMKPRGWodaexoh3WosgrlJgxhD9X4yFI3FN2
T0V/P+gVMq1uvL300g20ENbAkGo2t+Y3ZgmmIvbw8nZuI8gI8ocxtWCGrwKwaAeQ/lgptUhr67/M
/2Uprw0q2Hj/3yI10w+q/49r2DMuNhVsT1QY476fOAlX2OAkTHWfRJf+GuPuUXE7CQTYODqDlyoI
aVgsfX9/7Y1Dos1plHBSo4Vckeo7jwmmVFcr1ve79XqmM/ngSDdfwQEt2NKg7vxRmzed7msr1iDf
J4MREpMyDMQR8XT0dvKOKDhBjdTgUsln2dn+NEMvVhhv/rIfLw7hs1r3kEZqz32zQXHB3WRh8W1B
OquOnyWVIhzmqk7o9WhKQjEkMoYTpnX8sB2xfwA9rP/zzg4eEdMp9zajRoVqRwuypSou4OeZ4Nv0
W2F6FtYSjBtT4twRHCvxWWhI2S4xMzY0R31sE+Y9cuzdY8PLhfs9ZOJslilZMfAkxp96V4BGrEUA
gPcMKHaBfKAOuFauSGEISQB1aDlTHMbSSLUddK98ShFXytlRQ9DFdgIjGtLgD6d/eFi4Ie8sGXd3
+3yEffg6ESLnw1GKjmG2uaw3g+bnKafotMYhJA89XTBk+/x5ZSZ1dRCsMmc8Ru1mJkh6ulXb8tw2
TET6eKUssdpW/NoyHG2LxtRp5hesMxBts/Yhv/kfeNV3DykbjNaw0q1oepywokVCRhtYXgmthoL5
DPJ5nRHX0lVHjkVbtGcjeUTe+tphddXrn+pfKIVQTDewpfB5nGtM4587PvIvot7ZWKk0ZcOT95bZ
/L1y2Lr7kqJR6Pkg8EBDjlwyTtFi31lZcFAOum0YnTZPdDWux/uz6V0qlN7i/E89ZZ8ZKn6pLcqz
LoA+IqbxE2kBEhFbvlq8H+ng21tV1uaecEKDeC4SdO65QqCNRMs1IDIN0T96BUVY40BaSW5sCpZy
iGMNeLA1vHmtlZWTAigyqIg6Uo3GXQiJt5HDXnR6W/SdL/xv5j3Q/A6EcTX0M9LaAC3qo+EmTjgh
/fJWyhybwsvnbvE+y8ZYDihVDSgSuFQrXKS5yY9KjfPww/EFFodaXWEDZNlX+rbPNOUI31Beo+5R
s1Ihlsn9MLEeAFfJtAhHB/0nPAZa/Ub+QOzAVl4TU6lrOoeqPiAgCLoPE5na4bsydAJeorV2G4XX
Rrjg+VKRAV3DBltCAdZ+MgaCP/G5F67HFtKKO2dwjv1YCG61P/CFwd4I/n/+PMMy89JVtFc3Ayhj
1FU/dtI9nBXmeqkQ+nztIgzb8te+2+WU2AV6KmveMmfEMb0S8ogBXoRArh1APuUXdRgG/sGzcq9b
i5QlvfSCUEW+2JAkawVO3lHq00y90XJn4NI14IA2QG0M0NzxbEnHzfAD7bF8HqaHWdG5Hk18xZds
Tx5nlrJb2EkxURGW9kHi68HmYzyLRolsg7ClwHvOOn7sYZr6WaULSL7j+KrdjOJk2Hryv4sTzK+l
BiDKgmayneoSA+MnWjJIoO5xjy0jlNDHmbVyR3eOu7SZV/B3dK0uES1qUuD0TN/J4QCjJQdboYBn
OaTWns9aW1aKp50cN3h5CQUhjNy7xepvLgsfi6JZ9lOLvpN4QBQG8zVhjJXVdED4ZT7qYiC9rboO
lXvDdGJCiCAUzqZiQBKdyk5HGxATTmJDZuOzXPf1ugh+T31+Aly69Ntipyvk1TLiibs7UoBiknqy
Eaw0JQd3tSv1yUhRn1JuYJRa79ADeP8HsRALN4n2uoTHUNU15gSac0+9zo0COctVMNEqgUiNyKd+
074DqmPCxpmXeND/hW9Z3HBvAY0X9jL4JBrWxAMi/Fkv2h+PmM/IhyuuFwi78PNkqm74icuKNsBq
iGHLg9N54DlTsCYL4FI5zHsMAS8wSVGK4sOL1QU2fQbi9cJvDDw7ynV3uW0/mv4LVVg1UR4sKnHr
xNiIHt7urNgI/oXqBSdma7PXrLXVg/euILOQpP/0y+EbdBflA7FPwDFpIe8mtD7tPN0vwiE+4/Pp
N4n2pr7/oRzQ/6GbjvS3yks2iA1Qt/cWldITYui2t8cSazrh4WHhEmFBYOw7FA/BIBGI45i02h++
OHxq0012VdrqpWYIJoC8jMQHOmTU/vk9HD132iFAvpwaY+HG58iCkipTVVe99KERJQEXacJ/h3v9
J3fwxjpIhT82u5OTlpbPOir+dcc6M/AIcuU1F0p9/iaUdRB2t0eKZ/Rm84syLJaMrMq+TjHxXtAv
n/JvYWoxF0EXNs+UEds1zKLroTK8l6p7CE08lVHkBwv1BqegmzeEAq+E/aGRdLZccTQjldJGTcwb
nqXY2xj57sCGjyxwpTeTUrOzKx4Epzh92yWk3/6lKAb3UoQPDtUbbTMc22YWmm4Ujq55W8TJ1Bu5
6L/Lv1U3w4gvwfogcdjfLA/kHl6XSdjSkU14Rn836AE54S8xm8P9pOCP+8STXWBbZ0GV+hcbW9Qf
ev7G7rxBFGAG2eJG0fvivtL/iZViCeB82Ems7lZJxgsmUCymvdppioCt46ucSzjQqYN+QU5juAXx
p7rr+3tIEzHTWvO2gsEkl7lBwyZTOPvHhaYAG4CHofi8P1bA5RUboziJ7vgVm8qr8Nz8zbmmv0oy
vvSEtg/wZ+Ehf4HzzFw+5GZGWS4lx0hYbNLVnNCXFsOR7a30A2/oJ0YTX8ciA+xHev4gFJYMLmfn
M4tB0q1/xGo/njsiuRhq8yCgAqwCIfxvMSZavbppKFVuW2V1nQaZvJyof01RrR/5oJTi3/46Pb14
spAzrsvYRUuzxOXOCGUK1/2+2Xscevc1g1rnD5jXV8OIfu8cVc5TOfXyJZg9ocGoSQeKnZKZfM2w
SRXnliMmUr2rXH/Dxja2IFBv3Cys4TkMAKnjimmI7oClNcEjneWqXBW/dXYHvryvsi3RRdWYyWW0
pq7npfsGLfABlQpZsZAb7vlfV81FMJ3HssOH464T/ALcPfYO1yGDndWB1W8CIMOYcI+tU0pkM8Rf
Wfd2zoyOpAvcJuqGei1ONZgGCHhhkAg8fEW+Jp5VUO4VWmPopgkhjNLE9xLZfitwo6WjOev2PnVL
NVVsW7CWZtE7QlYCxrKCUPjNzr+0wj0JQty3rTuzCXHBFEF/ixZZQlyu+9Zv15pAVEuOPK0LMtDF
eoyF9PEe3hMO8ALYjFglW7zM8H4UEqcdROtdhA6RrDa3z75TxHyJkDgin2dzQN2SOMhpzcAc2h/O
HAXUaUHXOwA/dZJOPQ3QmM9hA4ffxm0GVtreqqvw4lB2/YfAt4MJRLiGRMZVCBUOR7mXNaSVzjEu
g8dSaSVFvcvYjBirkbKgfQ47kJKC2dMmC/LECPzNCRmFRXIFdn12CniEkFw9Ls1I5wvppdi/Zy5R
sl10ZtcMRAlYyPceOrLxMdRB62H965j69mrWwEBcPlkDva8ECq/IG/ZRy9QApq0j0lRG1uKqTb6u
u1EHBnofKsmhj9WBYbBhRODUgWw/qefb1gtoa2baSNoh0ojISymd77S8EWIJUn4mM7XRdRXx5/X5
BnRs/yhxopfMXLYEXymfO0dV814eEEq7rJs20GlkEw0/wnUclgsQGHCuVlFzmSlf1GNnFpT3Xw1r
WYcz7gs0j+0VVy91BzsqXhx6P0EyHOTRxpDaYimSS7CXO/OXfnqLKeNIVVPsuiXtBHfwNFuRGxLd
TeM1yKNmILn2X20dPkaXI8zfqYoOci9fGNtfyhMWb8jfhohKig0QyMOb3fcoY6El6AxLxoRZCWuI
3VSw3p7+Z/Q/YBdFq3sp4f0iEtWxkRwxMoVvvGYP0FNmUk0yd15aTkcjHn6+FDwYMKk+XhpmyC+S
XNFV86773dOm5Lm9gEHj217rgslZ/dfJv9aWY0zr5sO/b3JwBCKsAB7ajMUH/4QcTq8Cs1sRoCkZ
PtFougw6KVig/hUiG8Du/AOUcl3HFHla0ksAYLgYsbEeu83xuf1dAJWKdBf/FQ6EITk59HdByJh/
SZZwpAaIRJMZd5YaFuCAN9lclGz/Zr6MiggpEpxHi/qWf1kGjvFytbpX7PZ8PSTQ6DyKnwKdsJlq
E0//runVadFeBdEtTFNzjVsPSuNcIJ+gEiOdvOW77Av40TTjXpAw09CLjkoVtoq1jzoQ9dO54ITk
Tz8YKlCI92N/DladZpUFASG6eL8JdOLcvb0B+J5eO36LV3kSm/S13brG9l2vxDNBzxuKKkgosxzK
t8Caj9JmAcjUxKM4xsDg1qSyhBD7rFfLluh+bo/Zd78snknaanKoBygjRZ2O92Gy6RYo/7ppUhC3
3J5in9g9C8ko2m/zXZenahyMv1QFT3pYJvMeq/XKjWKycm11NEg1rKOHRnLvbDYygzGj9EcS0r+i
R53Ms652BvaSTn3SBKBgP6OADBmb9Z/Tdxhdow7aP6zPf+4H5Z5fm2o2HcdF4zYp6YkJN/LBYY3e
ivkdKkLnS5uBh/Fjh4d1GZon31ZSvbYK/F2Uq+ldBEOAWribe8yxOBI6TJ+pXP5HbH4nPK3+o1CO
tx+BToXCLLxCa/yizR6q+ghWcq1lQUIw0zzJ+YA/KNHmru2bYRthJMQDk+PFlBpU+3aLp1rDu6ix
+4OD6BZ1JhMxKkyWzTuB1prsconZmz6xt3sIBFvvU/o2zhGxNTEEC8k/sXOTmwpOjeDLncRFzXAz
hbFoZne+086Oan/C6hajWDNi+0elg5sGmNrTQajRY0NUwsZnVcve/KaSgRrxjGyxX3/7OgYVi7yI
jM7Kf6xv+mxD2rs5rm79unMhf9fsaoEILRE+CJyFyh4PUy939RuxOQdaHl4HBpDFaUcDFIzKMGva
2AnEXusY+75KKj+4ntp/zZhm+Fl2ULAMh+USQfxTNUHiybCi41BGY7qsqu2r4Z9RPrBeadctWlDx
nTQUuYz9U6cG4S8dhGDPzZyj2mMRrUr92ZvOLYpHBMmUlh948n35BmLTe5vW1p/+BDruibvq5/25
qzfwHksMCYuHfEu7BTo5XZ6We5lPgI7zd6BpbCInlTCvwiS7hNLwnCJkz9fepn3M3d8zlkedlABa
NRyMGBHYDY3rM8b17qviVTKM72noBVvdOin5ziHeJM8avrlG1iE718CaL8bcUBKj8I40Mb/dXTH/
HUuLd+B9lVc8H6R/1vthgGatXDmt7O7a5ZrFA7kZ2/QlMV7OkK8rP905y4cdS7jzDyljOhtyLC+X
xxIHJVAzDFaLRDr61UdpuPyFYl3/EbCoQP2eh3V5/Ei5kb1QC6mFo1Fa0m7SRW8pzKQsdpDTSu/h
9rTjJpShcgFugeYjU17jrZ3knLxjsKM2IFN7DHNTGvJwyYfjZRsRgp+q61ED2s8hdfz3W0F+rmn5
q+x5AtmlQXRXicDocZQz05d5Ck8zjZVUUKseFpqQalDZ3g/nWJDoBtO239NCG18vwlQZ5yRaPcMo
i/GB5FsaeVzyzyDtCQWi1K83BEbFNwHTHE5TpYcZd4S1cJgvLwxfqJF78qfL6tzIkzyyLUmNwtoZ
JoJW2JAF2mTfY7qBv+GjA+bi9CunoiG5R+/Z4Cc8jKlnBmBQLxbWfa42uVQU3TeLFBz+lCGJVGe1
HzZ9RyvmfiT8Ow9TkQcdpVjl2aUXHDrMskXx3PUqdp/L6+Y9aBM0zEetvu51t1fiut5BsExRi8lb
EljzZlv7WDnl7Xb35aZNe2CfOFxsOz9c5Ifao/SArNii2Bp4cQGcNtcwb7w4hVU7PLUS/0NnwoRA
YvugRpadQRLAbPK7ad3Wslh86aLMqHqSTrTGVlLy4vK+MgOvdm3qXknb+B8g7j9CFyQAkfbm2uxI
3H4GyQ8hNv0UFvnz0IJXzo/aNVaPrK856d85/XY8VMEQ4vx5yP6MAP22xNNr68GRmfi8OT0wofSI
Qik+TJLjY1qF4hehZve+ELFHJ4ccpWciUF7c28YHArvLZFnKVrSGPPCwT6sq/49t/tyddfvmgto+
560SwrzLc5v0b+6pVN+XknzqwLwJktAWLXPywCikRgVjnuWbqQBjc4b0Cvt9m2xMMOEaL8MYMVED
Po1EiqCiQAUeo3MMTijMEzJiWTsZZtECdc8y8SfvmuSLleNBqdaftB/oiQSsBdLdq/srjkcWVENy
D04i50awgvwghOtdJ5q3NMPjU22ZFOubqks2Q1S0Eu6ewG6IOuZatp0FLXajv6qKXw6enj5gf/Da
VeAbiCeTIUs7nL1v16tdrDR2I8u2An9RGxgW8Y6mBdtu+a7PtA3OceAAd5oQY8GpS+REypQC/k5X
HgQxgnQVP4CEYB9F/G2fo1+vB1iU5/85lUxbsnGBNr/WHczswXsXRZGNhUAuHj9zThRUrcj28uXX
nIZyGutSCBsBfP9LkB9rXZU4XYDeFBBcF3KU0Mrg5p37CuDEUjBQUfGOEuaBHHdItmgqBXH2MNPW
8FVfJCslYiwKBoXdoG/yqPNM/Hfy0DOoqp5p3tEMQm82Ek535eqM4riiQ8B0n0T/aJyaMwskVFAk
w4KnSapru3Kv9gxe1HGsQmWvy9sFw90xW6TrCVLM5dzHCpWjCEuuO3vRvHcUzM3rHr+k4C05jVb/
OZI9fnE73OcnfGXokyEdwltBDEHPXH9vT4u4/pH36k1ZFfcuuP0e43OCA0FfJR9pkK3DiQENbmXV
d2XPGNN8xv2UfPk3C8o6p4KuAiaKnXc8zim4JXDLH7ikkhavUOJJL4xY/nzk24t1G3U3dF8b/FkC
7HCVIbYqmzG73tHOTh1hjN/395g6nnz9po0QqUM9MFaiawOYInCD8E4cYobPelqGShXfUKRAWpHr
z/Yl6SNVef1n3ld/EzSF8VjpoXha0LspC28hGc04yckvEv7hzV2ZZyg2JLRMHpAH3SDpLRZU791Z
9LaYQ4S3oe76ciacgTv1KoTDEx2MlbgThbcU6OtKRrpLXnSa4uVz4WjuyKmLrs5N/3rXRX6orz3g
sX5Mqd/j4qQtYuhDog4v9W4YVPuaX7RPuqh6PHPTXdYzJuNIUuNL9/WICL8gHKGGsAKUAjabT/jn
eImduW+69xMNarbElqONEwUriatlJD5nxNqeUADqOJB+Ik9WBnCq/1Dtj4vXRqrnreh//Rv0X8PF
CjGvEGhGxgC8NBaTwZ1enFc1HxlpPsFy9lp390HinZcmof2XXmXagLnfiZUQsVCQFrr5bbZepbO5
cUBnm0gvzm1e4R5Nt1HQ1ci+h7ZU2EV5dJl8Ryf+TGweknMR59teylhmpYgPeFcJbVoXca8POG8L
fpUlSLpuwIf4W9JvjTi3wNCWhOJh1dB43xtRqTkmgmgEUHBHmJ0mvQWW7KuD7TH/fY3zLogABAwt
rahrl5MNd8jXzHDhuPfrI7TONhQdYuojXxrgjiT4vmR2bL9Z9EUyfhqHfVvL+MNMh/kjUzGDVmn2
dL/1BoLWQ5tGT9Y5dIjZ2gHNBgtbBj4aKpeC0rwG4V8aioHosW3b1KmXBZWHFyIzXBTltZ+TJJGZ
AgsjQEgX9LVq/b7ZOwLtVT63AcPEH3cjsYPo/mRrnsAwgCxJ0bu9qBHuHuMb+nD6K9L+d+4LXbiY
xfmYANugBym9kRldEXJTdAYIrT+NM1UA6ZxWjGDCthAGAhu/NSTPxiyL9p8eQIACALfU0SG5D7jH
B9KPCFLUUF2bWOvPCB9YoVuuMFF7XIm50JOk3MNneDjEuRdFXNOmrAp2Lf+by9dMxK9E9n0+LkNp
W4K81Mw4RZCFAQEBY3tiIRsuO7einuvlM/2hp4xpQFsSaMMVZgmF5GBUYcv0bTWdeAmbPXREeEd7
6ADNgqVINM8UNrcQPAN5v+pIvGPu8RLk6vv4cjSD07CXkGOT6XQ02VEHsMnYVTsDRYyIsvBa+dII
1I0INPCxzNQ8OigWUeSu/g2t6NuZX6We4FKNM2w+eZRi/GA5uhE3OqV1Tch9JiUlwZw1oV25Wrwg
WuB/r4Z7Ve1q30DHUun4DpwCBZPMS4cTW0cpDDBTDx21EEyxBnGuLMfYcVSN1gMz0QI/yU7pSTc2
Kgbn8b7RmU3KO3yxJ/rBh9LaLIl+HzXKmImdZ1iBZB86cpx0pwgUumwFkh6gSx6jMQmVuxkhfqpl
41zf5K2fkMSK/mScVwIYZjJHF39c+i/yFmWhoT8IwdkdV8Mv+oxk7Dhay4yhNKYPITVZ2TTLw+nj
PqG725uKYfaP5hO/86zOhy4ElJ1zBbqvJItFBtfCXb24Bzh8EgfJDfTPDbONaZp56wwnTOuGRRYy
wMiJIz9AdIFDjJY4T8TeQy+9I8JGh6t/BeMURnZ1/yuFdIyRV+Thwiny3Bxr/H/wp4NUwQsj3zQJ
YZlJ3Z47DFy2QSz4sEDX6YUk4zv4+djdSt629rH3Dq8qdIYkbED+19wiqBH8h3xpe3K6rgy9jFHQ
2kiO7CoftoamenDF3A+8phGWogHwcu8Adcc1c6/1pVBtrJgh7OB/RvkJf1Ca8i4t0Ld6bR1b9B2H
qYLOY5lwm4c3aLexOfbhmukWp20aP7VaBk2Hvd/G3tw6i4FeQmYubMaMZd/WIC0bfxtjoBidXG0U
0SvTUolqIiOsIe5rOLWzNq7I2Iw72i+KSL0LHczGhKWZwggDLz70FHi65U4pIje7/jWceHCdLuij
wO2kpz+bXnSm/6lWMjmhIQEWjMoRG8KugdyrMkjzSSXjaEwyV1RywfzVY1v91Ef9iTkae3jGwiNr
rbBw8nOg9l86X5zHWi6RIvKVsXK9+Jxb0ihXr/ErDiZxunjRIX5PF3wFsHCtSa3E821JWLcODkjb
9UD6CBHqMfPTNmBU2dTZTAgJxLxMEuJYO5HnuGx14K+00cw87BeoMzEeGVFwPzGk+v9Dha/wIkrg
U9cwtrVdcClYPLaFjKTFtTqxsgs+lNnYk14tYj9xRnVjCqI/CCQ4wLT9Y2sSrmlLn7oHTkiK8nzE
YFRdlOav9i5GKeL9E2BuJYlV4a4yRliBryO+WCmz1ANXTYhhhVYEQ5NaZSKBJoCiUp8Stj71v+mp
2XBYY3VsbmrkZCD0klOpp1E9TagDhtz0jwm9gprwCP3zYAc6PmuYsAOxqNPGsfa2iy/UKIzId41u
4Fs0uuqH9uZ9zJyqtsH986FBOM7+ENFFxHVFAUGnlELPfImNu5k0YWOO8N4NVSMEAnxOFBbuhhcc
ADSxchA5h06B4qqfQsm7SmKHjrd6NIAmYdYCdoVrJJhAjujBn/o6xhsLsuvlkQc6iEnDJMYEzXZJ
audZtLkwpNa0cdIEiRKZmH6oO7HqcRvH28ncfz50TZwMnefKZm/jZy+3tezAbZMRZeNBrHE8aFWy
eYAaonTNiz4KuQlsvZkBsMnnR+pEp1VdCapcNazKjhk+wMQini4Dv0+8Sex+4DmDTMRAcqcUG/0f
nyD43OPz7F6iHig8Sm1bm4WJmWtz04vtuZYF4gqnxu2HXCRmJuO03qLoK03Udcc4typGWTIGBn1s
kR30Gq9zbJEmdBggr0vhNn+2Amw/m1mlJw1Dv3+0XuVx07ZVhCS8IDjtV0tU1Yk6cfwPprpYRo6A
Vw22z78Vazswfk/Zr+pWjUBPQsVLz5/5H3fmeAPZzrWAuPj3EVGDPQWla55/kYE5q87Ifbslo983
b72kJH0qh3VmW8GIjt2wspXoizvo1ZgjKIpnkUBvOPRSxgl7BWJum0oQ6BDNv3ZKx6G3LXIV2BgR
WPWLBolBb1lAJQyItej+XDqq+IdUoEakOL/CPQhwVgJCCV9qtuhZrEjxaTomJjjMSvxecKBz+3Hr
ThgfoG0WfOYL2QpFkN65Ru2Emuu1GJgnkDjRzjXbswYnh9HdEdBCNkFaznuQwiYHZ+Yat52XEKsw
9+aHcE+bYH+pDu/3INwhHc7ateNdBeRZRL5gCrn2Q51IDm43k2ChMNevhteJFuudLOa1zMdUQDlS
mzazUJRo3HRq3lIxCfW84PLACgiR9g3P7CLj3bXQopQTNAP+CaklCsbzTVUmOre3H4gH09WetGRB
ub0OIZNMc+Ax6L2/Ge+nie4rSEOr1vrdhJMnMM3I8q3THR2jXEZTYo+Xxgv55hqJiYuVB4Fu4ks8
a8woSt2bge5eELz9zp3qDZ1+j1ZIdikg810sWkWj7vWa7dPQXkJavX0K/3XhvhCHzcPRzVwwunsj
d+tDu8C1tHnAVaTDVhaDetUbb9Ls4g7mFLaPAdetV9jlpnvjGMOObWNRuPjLO9gwS4LnOqGewJw8
3dZgBu2hARzMPu25YqQi68QOVzRp81IntGf5T1dPGLUCzjJ+Ec4VorLqJsrKoMReO1htia6KZi+X
x4xu9QnMux8GPhR9A33cmywdQAPEUsrrSbpYyymFBmCkhNYWTJNchrvnpNnav+mlcSFJsEmUEZui
dZ0k3C1etNNuSw+DwqMSpi18VdRk+1AfGAQ6MgKd/7wnLYBHT3fUj8GefnKHhVqPCU17BYbowlFr
2fIExIoefC6vCHnwrqMx7PDAVeRtCHs4WhNAS9KfVlB1SYOehqcOCaX6zbshf6a+ukaRAn8lCLfr
uKve75q8TejlwPDqgGEmwn0ga1GWR18fDb4AnqeZHeawRJrBd6Ml7bvMMxS8EvwTklGj3fOitaWd
49lSQ7r88PewXK1uBuKdP2Z8K5qPCUYX9YAaWcMTrVwcyiFm6Xn70LllBjPvb4ZaziWa6RhzCLaw
1vXq1qXngwK2wDu7kRpIVGOiw63682ieIiBpe6KONjS60L96mSO2+F20EGlOqRGV0xOZol9CftU6
VdagqDqcEaoL5wHPidDGc2A8Wv+aRHT+B8qBiGY7TOy8TPRayJsnnu/wymG0nU63+qMrc89x0gOj
QtCCpfyGm0laoX2WoyTczLL/WXlHYUs7pi/zNxs2HkItygdEjWPAZDbhh0OqdpMJrWhflK00vB2Q
K++ktQ6BW9ru4OGgH7wP6YAinF0q43TnUifST9IcaR2G+GHNN8OgyWBC8gUyuYzOafZatgZ4HtFs
UouWJ0b89n5Yxgd5cRsqLVVsAe0OG84Dsy15/P92gHEQWFRW4fUZoOKNJ34u4xQ55EFXy+xO+Iot
ZAVyTRM5neop3FFlBuDejazJ3vvONFhSmDvHb83vtUw5cF7Pa1SHW0/WC+gdWVAdnfakIrri/IrY
MPjD/XTZrR3FDIeGvA+sPGEOTTqGuuoAKIlaIQXRijZvRTOb11bCyrE7cH0pFsZBi1RNN/SrxcGm
nwNqfHNzJk8MPEf6ODRwNnNswRhZqEVtNPZlgzHxKklL3SZTGfR0HRBcfBNOAp5HzhYhAwibFIPT
b9oGFNfte8fyJelVsrKs418vFOEd8PLnD3ZGbtE9GpNfxNolxM0m91TI9ho9CL9ez8XiI7KBmsUv
jmnHsqpoeKynPlOSvn9VmFiibOawrS1QK85ObISjtQfqvOOk59E35m8LflsrACdYf2/g1tdtEr2i
F+BuiYw/FiaouEi5IKi600MxKk59UP+lgJt/qc2EwHyifCF4adx96z0YR5WO/aRLI4HL8NdBrQRg
nSsQMX4gA6PsZJ0/Hq5i4WQfq2y0ptE9Sg1P73KBBY7oKQv8ZGy1gaILgOtvq0NZOpxNUKnncRXz
AMqMkF2mMEMlaZdeQXNQo8zdREmFeGOSUPVoDBRWqd1tIFVNwXB9rbkYQg63svf6DiGpL24agoap
HZF867Ugt1+9F3DWlqYpxlz7l8Zi2Dh3PCKJgEYurGGDQAL+246n+cZy62PeYrt8QcQTHo4+RLLZ
bQz18WwSnob5KIgLQNLEUwJ9wfJuW3SDyFqOUZ7VHcCe9zD3Hu0ColxTZFdxPGSoZl/1EbnbL2B7
BqidB/Ar58nNhiNvqMp+N5ZRsb5+iArw3aRiPRfqsICJSOnieszwqT6IGhc7taMGjjkXAmYxwV1x
jUAv8QFsXqt8sBCw2Q/1Kdj8WsHBFSZ8lmPjURH7eqFM21bs3rEOUIRx+4631dvQAtgFLkAgkgel
QnEK4eJw10TXxUc+3JdBo/yfrfrQ7j6Dh9A/54CaFmyoV53N4sKaihtHx4meft9zUT1abJuke1y9
5CgWgksLUsjsIvdBBmZOiuAMTKz9o09l00c0JFdWs1zCwFO3kw1WuunCa8ee+wD8vsLfYthZvEVZ
Q5x6MckZ42xkSDbgsMTYr0OGgMZgYczDhIg/QZmkAV9p5IOSHG1LhWRjVnycos5AkCjU/xWCk/Q7
/ffDYd0HK0MdrPq4xJ+0Pj1fbTXhmk2VuR21rWbtsL98ADhBJ4+fuF06lFjJBZfrj4YDEahQBmNL
oyhzzQkK16ShwpLBh/LI/ESPVm3AdqqrOv6sImu8ocMLubhi2orOE5+wHE3A/FxduUjZBTvjeUsr
6dqsklAygLG14ZW86TocYDvm9nenzAUvbAmzvFSIZFCz8Nahc43UnS9cEdZK5w8GeMQsT7jdGTz6
y+fXWkALnmquP73SNTPUYaiONpd3Ekp6P8jEXmWX2uH7J1659cAiNnwNrqOk3h7tBOm68DwZre9W
/jCXw1Ys8ksJKQUXWIYaqcWlWJI2zTfDwF4giPzYwGKJAOykq+ocG+5pDdCDQvegOJIgq3opq5Qm
XOyjhV/LgfEl4PPyZPYt1pPBqQk2yx8WzzyD1x2tB3WNfyLV1EPHAhqnVvek7ZnEpn1ql06ns+Pl
iRxZNmE0v8ZcOTRzMXFm49yXuhMz55zDaIX3gEFZJ7neXp4rzDh8urK0em31pd0lq8ztiRLUhjt7
NXUUrMXKHIDOmq6y2misC2Fez6ihwPORTLt5w+4t8KlGUaGMSOCN7eDS17cvh14JcIDCPUsjn32v
uNcufDi+6A8TDx+7imduLCfTB+9Pf2964e77Hd1pq5e1dRrkEB+Q7wiy6KcmyuRQzw4feN8loeWT
izpC2z+ur3zpCzYJRR4cgidW9JjrPnDXEdbH4HRSrBAMBT9hraXvDRAcZ95QsGQNLbs9/t9JSDHR
O3HZjzuL5jxKCgUObDQIdGHJZrzfRcB/s6t9mcubXmPuimIqJPB6FsfhBz08yQ5LO0+p9JACK3Wk
KWGPIikFP/w4oWzltpxoVMzwinthjkZ5pM0AVmMC1hoYWJqMV6wm/QIO46nh2DYVvaw662IcUbS1
8oLNSW+kn+0tq0sIV6JL1Ig2GKaHIiJ2K3/ADm+4diAVt2WTM/TtzLQWJTnDLkPbq9dGhr1qNcL+
BCDtV5Bnrq77bb4WJGTBg/JdgByFshTZmfOxkK3tX5pW9FoDfX5xdIll8FbMBkL99pbf7U3ovCej
r/CogD3cJe3sfUt9EyLFV5G1b6Dd2aj8I4WB/SAQmpim1GiW6qyhgkViue9cNhi4iK/6VekdiRrK
xSv1Ot2+91GulFsbjbUfguCNL4dQZB2uNibpaMGsegQQl8uwWXRBUA7Xa1blosUbvWho+fhaVanT
ZOc/SKWWm91SAUgCvTpNPG/evdyRaaDH7Ampp2SoOftPJkpAkWU9ueIVF1E1SQwKgNsbKJaIgVI3
XH1TvUJGp03QELSkokoD8v4HcJAu4f8o+s1AjLtQrLXcIUeaZ3ODocG7Gj+YrHRbQe5dkUXZuJ+6
hWpvd9IHclJRlYLejXzi50dLsES8lJmFcbK8hV0pTZKaHYvsV2lnUqEU4s0xzcgwWnTGC0aeQ5BG
9ms5GBehFlyGRnO2xHhZuHkcxd40R7tcjaDan3z3H+/mhyy8b6zj/Bu4tVdnGYSWSDJkATmK8rxk
i7LTkDTaDrXTCtalea70A1tojTLMRDGkAWpYwQ1qbkfafM9w6RuNeFiKtQOiSCOHwanZYc8MCJdi
WKCJFp+ThP9jGlUgOBzlBdhFPoIJ3wIWmfvMNCJ46U+AyH3ldDn94og8le27KVyEjRfUF24zCHRn
p3it7xiQScDJYEvZVTXp9yXvQbR47XTVKJq4hmVz2uaArDSau4NnQ2M6BO967a/lWc4bov3NYi3G
AnKH5tUpPzuFgtfcdKhccXQhlhw+0AbvtdQgxjz/32ZZbwfkAWbPlu0EqGfKnOTxfK/Q8C6B/I5X
LTkSzBkYmld3pshIKUbB2Mb9hz1zXZ2df5sZMaIOe/F7MklH5mrs2zwQz9a7qhoJHr77O1SCEeqw
JAlGrvdy/AF0WARfzhY+BHWxO6vaLRFAa5YYMquJlJr42W+q1RJhDlH3NacVo3DI5pM+mGVCaSom
tWYNHZSs3hvKzOEacVALFMZRWXIu52W2CLiJYJ1Dt/6BW3lByOYSjKYUBg76lBKlyAZ8ux0JBvu6
/zi+8JtjKm1BUynrbmEufj+8Fia+1301Bc/t6wVgQAO8zpZkDIUCK49blb5izVy1hTH9AsOjAAKy
nFLQDmS/nqcgT24UxX7o5/hOz2iTB6JQ9PcaF3OT+TcTTilz4X1L7AX9D9iNzakxf0Sxw377b6wh
o7+DeqYcJRUdkwUFQzTeENl7Yh1asByl5ycXvC+RYtt2VCYExpKyzfRT6/Irp3jJD0fkXas0/S9q
k/ojGWDV6JHe4rTV/WREX8y76p2F5bR9N88o6afymz4xqZXCgdjQvV+thxIAU9EFagdZ4m5qpvBm
ejvx27DKERCNHLgH7gr5zRus1Kl0TpFMG8dzVv2402bUF2eXDaAxQ8vyoX+mEvAfmXg+dZzDRXLn
4EanUZTI3zm3ye2GZ7EJlWwYoQCBgE1CuXwRxSZvBZWPKG3zs8rKG5Nkd9YKSchTau3MhUh2cNIx
M65lSqCrQ+TAjpx2qbDZ7rBXnk1t4MRXwQGPYnYvKz/m50PWHRwavoE2tFYWWQTjbMaj0DyEQ2y9
q3c0MVZf2abkKLoTAZmRSSc1EgUnItnoDSfhs8GQTZwnLrUF9JrYBUAB4QETmwxBIVN4U4+5JGiS
jLBpS2GlfYbYpptIYj1xSgnhwejkZ5fs2G8BiucDUic+bOyiZvdqVZ6gx4pj63zDWqejNCmy+Kdk
GC7ztZchBIssRG23PF3vrpe40le8yvsAR5JpzgLwQ47tNgOLT09liSQM+2rkY7Wp+oFtA65jZ+r1
XqTwjfalPsUAc0AZWcodIrmPST4nqRPTEHSMYw29cMPFi4SvEYURRoqeTrUyJj/fZr9Ybv+VzsFf
ncDIRy6qRRGzAeNyrfhQB44QXoMT3y/CQi2KEnlKdW3x7JiuKcFK3EY7NPxzQpK9qXGVum/89hR8
tpmx/UDGM1m9ifDNRq/dCdDTSt856txzxd1ndpjIrIa1iGz0wwWiYRSICfvxEDqiN0NRIh11cRQs
kxmvaEipJoQbo4+KdgT6QojtIBl+WBNWuwkHRGe/ApTkUm4YCN3ZMt8fPTzujzpRxhurXpxI4Bb3
IVAcV0dFgTBNjk4MU58rWiiWeYtEWSHJwy2I2P2NJckePhJLLVaNOkRdGNuMtdNN09iXT06aYnXx
B05K9hzom/SR7E9O7F3rMbiibfVlj7eGgjPKJHWF+8NllvrsYPAng6ucn3MW0L9ymgAmbxJpcwWs
46eY32ExJS3WP9UVrNdK8wjfOzJe4XJcm3q6VQzkGjSGw/AV44jKl8o4poJH3Jce81lYFvHDblKN
JPh3gsrcZtVjRNmDfoq5lNCXHRgH9ig0VIkExGVOTmLPjPDc+Hlm1ZwCsexY2dE8ySdJmCFs8dm4
CmcbLZZShAQyfISMm3hbvqy+HFyLOKJ6g02y+Elz1zqxLAaq//BWhO4+mu9P2KA34J87x8ccvFAV
Wb5GrhtlZZ359E6l8wPFDhiZ5YGpGKxvXp5ni/LDxyorMVhLxSYyDPntTB22hcSQyGH9tpTH5Ftf
2QcCIkOOY/bHlq25UN9rfVx6HphJXBEEne6lsfutf1FCfTl63bs+5HG0xrzqPLE7An3wAOB/G5gh
+0fM8pJ7xq4lVjvBKYdA8/mzjzVMIAKbCghmnM8TE1vcpmQJzanS1aLkOlu53dBYSovRzHooQ24D
zWLhj02JgtK541AH22fh4gwot5gqaRyo2mM++TPx2TM60EyYbhwuDj/dHFo5lQazd7k2J42JcNdU
Mg99SuG43GTFjPuEO8PNO3GuVhVkX1GG6NeTLi24fSLe1IWAGnHjD7mjeXPW9kZ7IbS7FSrDuBzb
Xo1qb/YyQ2acMWEpMF3pzWSVBpqb8DdQysX6i4IDO1EjyB2IHmF9r/wvyghgl9y1P60bxUbzTfN3
IvNsFUawStBH09PH4KO/g8flCEW3N81q9zu6yf6ZnlqAgpEsZaUvdQxhkerutLxQuNdedi4RUMqH
OlVHKFoVi7Tpo2xeaZF+MoHoqxLBdskDPtz16dYUtZ5sOQt6/GDg/8yyE4ggjt0hh3U+gEaDFeLE
RBbybeUquICnam+kb029gNxDctcyrrBz6sg/GwT5sp8Y7lDhROdilxjWkOtXZrFeAN2olCrm4mD6
UR0tcZfWweXGcPlafAtYhh77mg9OcrrTDgVUceKjI7e131pXMDdnvAWhrKhKdYF+IP3ezdQlblTs
o5AuejH+3AKzrGrXz8jyjgrH2Y53zTNLc2IpWr7e/QXva6apCM2ma6YLS8CODwI3JPpxHUae9YDQ
fb5HZbY5EHzUjyTbf4k1qKrsrOcgL5ZXILOOWpuY29oscB2bYu2DntJD0I73qR0ko97lGuxF4TFJ
ThjVqvUfcOsAQyHiqvWUeJmx7nJWUXPnLtpj3FocLVkACSEn+QF6G6WMEbH4uqP2ZTyF8GI4doz0
HjKhVXycuDv3wKAW6pmg7RTldUKCU7QaIwWLW1b0NtRC9rqqA1a4KJJ1IXwugehMjOmFor32Je/8
fG4gYDsUbkzy4Aegm2GFN6WyPmNR3+N0NjTfQd9pDxDp1D8MZo6uhJNFQ0LRsNQ1D9BuKYKN0hYQ
u6rHwlytuRnLRHXKcYEg+NQ6OOnHH8rWzn89PN9BCtKJMAxnK2EEM0QLpUD8HCudWCqyP7ps6u76
xMgQaxfZUGYAVgbuVTaiOwwm2CMfXTEHoB2lOpH3xw1mkRueld0pY7WlFP2tTAzCz0WqW3b6LFZ2
HHbtzIcrj+81aNvJJw4AbXvpY1q754nyX0B2GIrumkdqHESIMgKelxTp6iw8VKgGSru90ZrewSSe
WepKfM9WyOQW6eYc2TNvnkEfkTwY4alLIbOlYURR6G2PbCvFA4mC/5nj/W1nI2aD95ThQYHCYWi7
5oJ/ch1GoeQOtvvWkCLMUsIM5tcfQZuV33mhDANJVeensBKlfbvnISBRHgLWYMo5C/DN+njlxQ7P
vB6d+VjjKuoFsu+VGVkJac2713LACZk3Nezjcb81/yx+2S+ZBeLrlNh4jmKBPqPDez8FawoA5vum
tSGnnmUbyc5ObgzHIYFMZxgzKz18sRH3vQr+5A3dc5C8rsqkFonx85BmkmbpiZK8WD9L9UoMWmKC
m89PtY1GPhyWwOYiB7JpbYFqE7ZisgG32pp9051E9mk1h0QrMeZgw06Sypt1haos6o0QkeZKIYFW
rsVvuvMtgPZc7RP6FaAsX1i8ROJJNr4DrkNSbX/RjJ0zWePqyD91MPGy+2vYSfrCTPDZzsoJHkoP
sv03g8COonLQX0uqiCcPbH7540R/yoKBYoVGO5FEQD24dnTI+t6N6m8WX127fiysSXuWrxU7dOVk
o4qbSJtMFqxPakNuXfGrVx/gOzAm62TQpjJqf+/+197jivdL2HDKd4Ff3Q7cP0zrPlkg6S6qTSsv
fJc1BaC5hYnmAgNmKJPKCq0QwZoK7VZHGvyyFz9qfRK3WLD6sblRiP1/zvklhJTzA34FLk2nsnZy
VRU2fuT92Eq5PSORCKpH58nyezncCZPqkFnN0aEOxaMyO1iRl79JBomiXKUZ61HdMLfTJ19p3JFK
9/asDV8N1vQnpx8sUrMNksRwu1VeA6LybRFqslzJWnuuSJOTMn9D1OrDTsRf9MkPK0vJFJE0UouI
ZFtpLaH/KEhFQK51alGzPedn3bWIxHCDwnDM5lpwGIAgod9c5cOL3yRtvmDrIMvpUz6fMwoRNkos
zYyYvJhJIlBKuIuUbTZ3cIZkteOW9V0U3J/UdYn2eCJO0MJ22prZqhWnwEADPypcvCMqdCjMyUqM
hwoeaUv918ZoWJ7SdCLSizLWq9Bid12mfwg76lwUSWF1ahHEN7AQJNTAwfOXJZwK5tYrRm5+jqFg
phI8y0r68z/g5rstY0VL12O84ao6G8lL5UuQ5G/sDAQabpIcG5VEatqsrmFTKAEJUMXITGaToRCv
ri7Pxn9PfcpgJfYpFoVDYvtPSkb4nJrN9eT7AdLGz3M+TYka8HNjqCTmjXOo0QD3PjwqLpM6GhDw
PAEeAA2nlHIQ0596B5W31SmPOMNBiKSkooV6OCWYLYghBffMqj0YUho0jbYh8/viqO0i0e4yncqA
CM5udCE1d6+If5GPgHSfhBB4gsaIxNflida3EmJJVS605zhfBSfgMXP518gv4roQ5TuLT9YsGuNO
eXizA+twRANX8FTZyjUwYATemmuEgpnnkqohuRtMlPp67QiU3e9Ps5UO6HHxBctm/mfnJA6DGldo
84h0rUNlXgmkonewJYZuH8dXJ0vGTb5FBG2qxMq6y9BPgLcUAKk3lKPfV7lb14SrRYCAXmyFM2L4
NFAwZIubFTNAq205VS7W7a6ujVNZ7vBf7sKsNIc2+REBUf8A94yC98FGeB6hES2PVl/zdwbUFWSY
o0StUV383qr0KsHJrPN7OdTQvMpecrhF0G1oNm/K2CbLELCeoyr1PWJQJPp9TwWL8OQnIJllex2+
1RtJd0ht7nSCj3Cl4Rrhgtb1ZzVzC05i23B90s9GevJaER9JJ3vK5CVskNhbKlnVrsY/nWXzK4Rn
3//T7eeCkUDv3apJz2DFNHK33w2m8nt6ahX6AcHdnIj6coqQF5BKrgOMXq/TRvZ5KVg4/A7tIEUr
ni7lglvI6pbe5AmHIIjxWUAJS3QuG4Y301zdfsV21oEG5LvkgLwZ7mbTz7ZTIbqJohGFZKzm5kFA
s+/xjLhXIgzgDGDHH7mn4aFRSK8FjAghsH7+5sZv+/sn97L8m2AFc0OfLkus8TLTj1fTNHr8ob8t
sMqqOJgJuDHGMzSc+naL8w75aDExZCE7yPehh36kutk0ZUxD6fMdhk7dYrtpI/ejBqH6mNaUHZ1N
3ZHQzkIi9NbU1+gWijvSZgchsXo+1aFMaII290KdAiwuScRc6Lpgz4MxOHcACDpF9lOl+HzoUFuG
hZzqX9qLnm8mfFss8icR1aUgM8iZlznwlHONmmTEtseA4wH4HNQpL23jsnEL2Sfp7X+WAHIStKVa
t/LuXB6+dEXuV4KUDnloNPdAHz6I1otQt6qlBsT5yrxVpLG0f+qk2qeg1iRSALRjMWO0SX/eMfaw
tVWSx7W0GtXvRV5BLSfMb9/eLmmPYAhI5lE8QCSR6HGkkoYnZcKXpLXhhvgoGpgfOn+SqHg8r1fw
Zn/1TwY/HJv8AOwLQc/6LjlK3C/4/1n4i1rgKz0/Bi4JO8HRPkuJKvg4VHJ80WEJtcoNsdmfXpU0
5WsRnpJ3hsHGMeETn5islVDVVeUlW2AiZiiz+z0SvftEfNZls7+AwquJLz3BwkFNlyPKBO3FzkE+
zDjTUhFgp1oNZFfCkqa8TqD+lFrwSP5JK777Hd9325l/kJ0SzuypHgLsi1MgECz2IEUbtGPVJmd7
3MRFQILC8gExDv3QqabR3xOTJFt1806dX90PWXEFlOiL+XSDAT1M4+7YPaFl0B2cB4cdaLRiihyj
G4UrwO5wYKXWn4VfygfP+mVmqo924R6POQPvah94r2M9dz2gPlPdGd1TIlMV86usQQsFvfJGud2Z
zKL0mgfj19bFtIT2hfmFPA1L1Rqke6GlzKYlyRhl+Z9nN6NLXEeCmmx3vCaslYp832E/UKjeO4mY
qL8jWQxkJ3OsLE4W+MD5V0ruqz2vjobEaLeIG7q4tynsF5Mgue+3+BM5cGPM7nWT6xZq/mEWihaI
WDKylN+FzOB0Vf4F9c9QyDktXxQud0Kkr44p2U3RAnLh+DzCTotvJRYFps7uNLbbXiQIUqQJ1Ix0
c2n+/mFWu+7WYiRu1NmV7FQpnBy4cn2IFD5fujCA+a/fqw8gs/0YFWqW0dZjGVI9aPXwle1Qd50b
+wJAdMj+QJFc2k8QN46XNPVMwmTKIUqqHD8SBw/x4EmnhYJt/7YZioAVPRFMSq4t16uJE7Kw6RXP
LUwERXo2t8sKoQfQNcQwd3KwpVQlmLhO1L08nKTWepHN6PiJUU2vaq+FHz8dfslpjKRM0pG/Th4i
IzzBLyPr0m8AyolcIUY4PW8ELBCXk5Gn48V+b9+NtheK/vCov29mSpCkdZjd2idFzjN/oeb6ivqN
w+YBFBBkqZCnKiINuCp1SSWqlLPfEXsLGH+a5KgmsshBfZbr+I4S2SYYOp72lGFN2EgCi8Uh+6qV
a0JLuS0O6SWZ9JfaETpdn9/EBXH+42yxAieDxqQ7x9//kKIYBFTO2b16rK100tqL31CcRqEga38P
TML53fPm6a4EQNMd2XLc6gbG1nkX2atgfg6diuDitJzfa/kKhQtKzAJzzM/w4mLAConH7EtLFIYp
mmmtRJdz+/QZDUWiwpJV+T2T2U61W8Tj5m09e0DjkvZyjz3jnTt/fBPuDvHCtGcdNXcjU7rAuqt8
WJ/3dlvqw+3r7+wU6r1/M09CcfLU6TLIjbEoUbc4FdnOTcyrx6Mv5hsdZaJuEtHlTPCZTsSELbZx
29BcmRgc46OPJAR+jaBPH1aO1qCM6q48IGxX2NBAFnFUw0iiyH5DcDSlcWa5VcfVd3ASQnwjXrRd
VFSy7euteI1fsQquhOypQzksv2uL7uAs4HPH6x0aU4I0FbtCLP6ZLzH5dDnWS8lhv2fKAnHsBjCm
nhQLfeTV0fYkSRtYURI1lJE25Qd1ofQHBArqzGKmzUIp0aA+YNTpdLM49nTYLNqri3MnRA0haRuA
Crdc43Wd9W9xH7Veuoy9mxYUhF1HPPYIk3tCUq0zESXL57GtVP/1MMByWCaGLQ0au8wepTVeptd2
zJ8VfHzVwAJj0xHtQ9XqbODswNSgLRambwAwvwNUdGJ2+AeGsDZOcCfKRSXT5Ax7XP0x4RWkT2J+
NOJknYSSu9bkKOKW5zxSYx7H1zgyO9zKk+CoOINZqkEWCTQ6hoJQJOfi5fJd8QcnXbt4QbDepVRJ
lbJHTq3tvT4J82EmH0rk80vVLZ8Qk3Lf3AvV//AG5ynTaxcYyKfjKL6y0kd9R5LhGEjHhdZ+v0F0
T2HSLbl2o0zuVbJcrfHx4AHzDgWXLFNvFkGuFIb5gWpoUt8Rn1wliHLxewA9FFt6m5y/pTQSNcec
7Kf0RpDjeE4ZRtuR6s3nNW8LsPJWOXQjgnTBMLwI3du7KzTP4bfHupI45yTReK07e3Fy7CBQHC6K
aLdJOSFODIR/nZf1TVcq15aoC/pnA+fdV6lFKtbtSgSMSKWJKZ7KpffkE9k6elgVIxkCn1tIhPXA
guQ1/TdSTQnWUf79Krd6gOuvmL++oI7i8+UQTgOdc751L8Vc0NRVyL2gqueRGFxIlro4c7td0Ejr
lWvYJR5j51DMQBk88odMpIfbnEa8AGrrD7fIwCX548fBNLDNNTIa23/Y8tTjA+yXAXKS93dj2CHO
jFB1fnxCNBdssJpQC94c4lV0U98T9O5TLF92rbFTgSDHUEsIkcHtcI5WpR8YjTpjd/gC+Ni2REwR
MiZxTWaLwh64jBgcwHqg9+iezZDEZgJtPkmFJNe5Lme5WcXcTGq9pFwphZcLBaRqHqC12soZ5Gqn
18EhKAM6tkA8LHblghFE0EBnVnozGgijqEkiBXqdrkD3xhr+eJFjK0qyLm5P/O/vEoIfHCkVJ2Yg
5/GkwAlqtNgRULXaR9+2Nxd/XYTsRd1/8kKQ8l8CvUSV+cN7KPbu8Z8Iut/Mr+raGm5Ikz8p9L2o
gZbmHzyQWAqgPRoAXMd7ufVJJJuL+qj/9rryfYAbPlvEabtEQyWnSnqsBBOUMnI4VyCWfnH8aKd9
dTOre7R3GL72XT1Xl5bAuT/KjS4YwsY2KN3xSySYesHT3IFlT7gKqHqCBgMD1/Zvq5u9WclTrXXV
liSGtKV+jGnxSxReHAMbqyL0bf7w7aNXJm3T0sMwrrrewFCYKDQBC/AF22slJ22Bg7Ba9QJ52vjX
jFdfxlTi9mRmQR+Vfqpc3XDYOgx5S/v+wuhI+pHuiSGMh64aBsAhQ/YRwkHX+te8NJbJHVIb5Veg
eCU2lgnQV3S1MdCMFzv+cZNQCDCgLXkZUIwYr4GMKdw/Gpjnt7xdyV6PkbGM/w4yhow1UrxgHqEj
CJ7k3mK5+uWKRtsWXyJmGz+xHG+4z8bPNWDOQkKb7r87XK8z6lRs2rSl7ZlOJhalGatZniH6zGFu
hb7lCCuBrtIZAGDAU3k1r3H6pjhPdxgiQWun1IXZvGgH0Djr93ter0yqv7tQDZe5isO/I1cTcduB
hjf4cKxfPW50Xlerof828bSesP6WF7NHeFOtQWrbAw2z715WxTNqDTuEA6TpXGMDMvpJc1Ufk7/a
b4R27eWlGzOkInqOVeHXNKPLYBf8cdytEfwRih/0zFojaKPwYwyTM0VGz3ttOX1q5uwPxzhuKE2C
p/xuZmwWreLOMx1cv8yn8RvLg5LzNOrlCvk2AW6NCA4JOA5htrshBZe4qPh0pZWyoDdcLCC6ICHw
Mg6IorB3122D88YxTe2vO/3VGZ7l/b7Qr+KOgRWytoW3rGi+Sj2P0fDZkyI1QJ843gSMrDfgU6Df
FSWjZWRZwV1YQqZ7akSa2SRsUkDRj2pcoCiEJMORd9criFdfNEtA/UZ7RVgYUEKtaRF9Vx6Iep0b
HoWECmPeEk9UoBbd+NX4qNN6lHjuCiOaTCF1lZicF/AKsttyci8cl+ClH5AtSKtazeLsmGD3RJQ0
5Km1VCoIngT4EtTxLhRfpTRSEmhw9wN+UGgW2giz33nj8SPYDWQk1ejH2omyqBh86nJW3QnL6V9b
eI262V+gGcjHmRmRe50p90Qa1Fq/koSqDoYJLYftANJiM5anpm4fkrw+xzLskm1Z2li82tgNSjgS
Fs20l2UERCf/JaSDSJwU1fms1Bj59jygE57OOC98DWrkgNkdOxpehRlSL7l/HNQmE3O94xLxrtsl
8WxyycuAJ8H5M92dG1hj1U9nYcOYuSzuf1LcPVMtGqWa6GOLJ0g+VBv0wldxbQ+IZaFbJQbL+cHN
VNiFArvV44gKihyNua2nsxrfCyoTqvemB7uGsrpFLHKXl6F7TLUyeG45BX6RNUeBQg8PIco+SiMh
o7u0WURcN4ubZHrje+Mcw6H4FvN4QqOyojtcN1uY9/sQphWZ+Etf6AsfbJBcm1sQEK6O/C8oxEYY
sxBFD2Z/XqE5dTMRQbFMlmKkBdYWjtRjhCwsqohBv32ml+zj+p5bVL7nFfz1ckA94uIECFuNKkNR
rjlWuFoAEKJSwS7tpLh23eMRSo18Rj5aHIkeJvGWW1TMtpE07LqrrNdVSg58CIolmkBREfGRyLOU
9w/ykCxbsOWubOH0ZXUrqnvHnJbRKpGlOqkAzK4e2HEOtlA94WPF4F38DWVN9V1zdWlwp/MXSUTe
BgQfYPOGNnFOmKk6lYc/FSG4SxrQu5zT6NJxqjFewEL/l7Vx6YjUchQnPTKmKqPMGLpeJlbpTU3b
JPWuQiuE41Gjn0GTLtcbrzLbieswazn1zFka5TQF0Wr51RRM1A+oQhpVcj/LD2xuA0ddsZV5JFke
Y1qr3rbWwNLkksIq0p7R7R7HxXWGXrqLYzBe3RYauTIsyAgEUtsc9R+uQug7dMI4QlWMOC8hfqZ7
eY6uqi5pXUFvbOT23NTZ2pzcIkADsTVUpMaASnhzJU5JG1uruVvLzUN/ZDhCqO5GroDkwDw3O7ER
y4qNaRXbkph44Vq9mZAfQ7rzjNgXuRlsFB0UyRMBZVtaMYj5zWVzxJIQPTU5M7DJD8KKNA1e6eWZ
KDtdqSQhhYV1wxM7tkBWFk8D1gFPvMUZvOqAsmojaiUBAKfg1pt5+Tiaot52fmPcu91uo0kbPfa9
wuP8807WvrXA2ZI7hE6zIfKACfMGfT7NqZIO81OOxIFCF7ah+YW4zZABQIpkAyOZ18rQsU2tXzGn
Vy9zoi67MAyEvpAvVPuaCVbUfnlvHD/L7NFl6rLwBKB558VuFaE0RM8NDWeuUk94MicDXcxjU3Nu
s8SHfpehPFnAIM5fTHRrK4ABaPVSAjgQJ7ExPHloy9ilG+hqpD5rrePjU2ShqGNi+suDQvE/SJLu
GGcVcOxrLWxUfVQS6r1cPMHtv8G2We5x8S+SIAz6GF8AgxQUMa2O4RIliTiPSFvKu3kMHFNRv0Bo
6lwfitoXy0II7y3KktzpENVmh6TlzzZs/jLYe2Y2U+rOiE6so4Ywj7sZ+W7giqX1y9N/c4oQyjqT
CrKj0NnlDd4GPogWAvxyaG+FZA01OmD5PJv9YNmpOKdK7ds/rrc1QtkJTED9isPUrg/vuy9mg23f
lGvbNISq21I4cW51Iwyhd9B8n8W8sSxqrrAaRXFwtZx+ZNCUhuprRLHauKnVfA4wCqvdwm4pdMMU
dLHcCzh7kTz8lEMixxeDGesA1Zni9JLi3H94gS7CIam8N0GYQv17dPBVgelCL3KFecYASNPiRF7X
NBUosvqLVO7pccWDravbW2G/hLNCDYDVzbNT4bjsmieNMGgpR6R12AlAh12Ij+IxOeRVPZq90+ye
sxoLrQPbq6PtykuHmgmdGjXdruw2JZjyjFVG3UgI57reTABYaero4NpZB0pgZY02V8mMA459tfGj
3dSsl92yWaqSk22WfO/YMjUORyOFTlNtfKzIL/q6Et1Pbmi9VUgtnTGVW2JtNZiagRtQtDqchKp+
NRillZqNK75ZU6rmq3X+F4KVXOVKBk/FDgx/tW/r2vw6A7FzQy6itY0eOl0y6aIwYPGKguwqFv3C
emPMBRrcdI6Pxz1KzKtP077tb8cRmX0qDxX6gh9S17hy8T9y/23WcSAcIcsB7qVybLON2Fd896tN
owaxHNui/JoJgYfk5B8FTdTbadPOIlSYDKMwXKBO1FTw4MGGoHJjXV8JJZN5f7dqeP0HAg89Ohlg
dTeoFm950aun/RQIfzdjqMwwjq2tZMxM/MUeUoBHW3W0zx7O8NPivgoRCFwJW9mdT0ukJP2xeJnB
XeA9ZJo2nZjV5D6nL+CMmH+4OtRK+qJ3NiCyEcHPySEP9PtiX5AlWT90/Z7CqPe5uUdKZM1EdJUJ
P5lZOLqIZQ7svhnhfNpEV4ZXJ2CFO3vmxCVq8E9A0YgwMbH9PoYawDi8sHYRTrucm6gOCrO+ab/8
OzHhL8Ttn6lfi64i0ucbC/ftdINq7tuzUXgqWHb0suVe0jxCTGkqZ32N1CUJzZfT0qJMAB41qHmw
b/W1LRhDLM/CnarPm7ZQEZ2ZublcxqGE4vCW9LUqgb4WAWZbrTgoctkbPDXuz0QVXnXfhoDtLbKM
KWCQgSSbPjPBmLm1+Pb3XYFTWibbnDZ6qq0pBEhA6at6KuR52Y53GQfW6dIi7YRpcywHGUkCqEKi
koGxX02I6em1TZfK7Gv1DGIY1Jj1zDrOGYP8Wnt2nbjlRFPAafqzVVvRx9SsPdUe9SP0X8nyIWev
bkECRyDUQQStCrvjzq1sFqxM2aD4CiqXqEk59izPTjy/w19hElWuHOk+gX1rCl1qY4/I30DBOerx
5WTCyKBQzkZK2DxrvHaETVKjAf4WQIgGCD17YxV/bgvSIu9aRYlOgvbarx6Fp84BluWFh4vQeATj
2j9IcyxTASZ9zkqOgWrcMcqwXG2MpWCQfLefTyWhczn0zzCTR3vVFSqUnNBOwvVd7mSE8Uwx36la
fEaKtpfwi1+bhveTSIylMSZjRnVa1HdacZzoIxWjknYIWzEQW8j8r257ho5rnPPogNdODGCwvrff
SkhKyXwKEm8vX3ELaEAw45S5RBH8x5ryqVvL8xn3wHybGr8puXcmmfKsJeCoqjXdZ5hvYuueI4lv
xhvq8HL1a85rau4pfaj9Ghp1b4ojOaj4mtHvMlANX9VG3qslYcw1hqt5Fq3WqR1Hxgxv7e6MsFMM
hd31DmokwbwkAAvXCr2Qhl0zrDtvevZ1n+teH+VRJ9XlevdXX1hyRXHueJhHhpekQTTU4PWXZkY9
2C5jAj27mM5/A+lsO2p5at0U4yOUr/XyXzO3Bi/BG6SlK7wxGbARF/GAh3gy3lallFBPZCFDwxA7
KQtC9BxojYcdV8y5ZRw/7NCEop3ftVVnJt9O4E0Kars8RftNwtGq9pswrCuFq/KREvgoZmYlj6OV
lebEbRgeC55vnRAvZ538r4OUyyMLbvG9r8dDIUqf7tFtiQnJdYxtO3EicS9pcfol+Xf+hFaZb+kE
OPGFsgRdKgdPm1QQ0nlYHHiuUzemGSUq2wEYxKaSWzS5vPVpgd4FiSwkdTP6D4BhgzjpD+XcGD9Y
5rM0rktuD+tL7qQ1o476nZd3UGtdGzBFHZm54DgVQdFFOKnLDIW7blx6yQGtMxLwy1ad4SHLYtZG
iulRgtLAEOWIMY468tTjKzV/uq1/8jEOp9V/94K6+jXb34ltwFgsTrbQpBmZxjNqtAN9aaaDyUt6
SlcKSbOc/nQpFrHBgeX1NqKIiczIBtKSIuZPrFWgd3S6wZrcGND8eodNNj2pcqjNV83OIv8tkrvy
A5Ob8UeRcp6yREZt5QIR8gbNYJQrOZN7nROkO+UtZPQnp2rPPOO7PgNcfjgDDxk87EG7RvkdQ2Iq
h30yhbqrfHj3LRAngXoEyx8Bsk8Sw1e2bK3vH15HvxsH026P11KMYhh/kpkcBfA4eYZCiL77r/WO
lFVeIq1T3GBiXkoh7IZ6Cjww7fCQvT56lzwR2nuk7ZacOea/cofZCbuXZBYaBYR9C3NJl3L/Sy0s
+e+ALEFML5kG+qtp9fEcSmY4TrNHljDTPhjSLG5C8OxDldX9orP9qgVyCxndXaFDJkzK/UyuHkmK
oUcE4ud49k1p9oaRkiA4mdNoTQzrarT7VeX+IJwDP7TRX7ETsckXv8Q1yx3ICb5Hd50YsDPrXDpv
kC+3q0wzGso6hsig/6G3sIMISSAP1Wq45lirTjW8z1Z2WEO/s1gA21aL+HVDttQi9fR82cCgZegJ
9jjvtr8ro9aiefUC1K9ObrHCeaZkh8+i9rkNtew1HGdIdwJ+0/4X4iNsZP8BsUT5+lp7KlPI+zf4
yc842YfI3gwD2Go0CshQCx/gBm15ZZlfZnsXM5Oo0xxiWTNzMsjS41fqWYY+uLBQm8mraA6SHLgI
GokDd4DlJTdfMDkoca+JPKIYGoN+4m+h8J/Gh5WWIVTx9Z+uHow7gveHvhI9mXCF/qnqtct6ZICr
OKSstK4o8tZjZkkTU9jEa3QR0mck7hnWl5IiqjfW21luQjWk+onswqxdwTet1fQCr02t70TOiv9S
QGMeFWCoiMP7kuqO73r84Duk0bRnmvmE1h0NMavcBU8nWS5W5oXY2AVlUI9U9Q+Bk29reQv7Ee+K
TLHH1xEz2lts0FArpaxQ+1mXzc23gFg++IokX9727iT1QE6r4gjDlHdguJzxCoU4BE+elWdAqBS7
SxyGbs9PvZicdngujWBIJ6RTgzpztYW1CIJH72fo1VSjpeeFRwsh9N9yOMt5rWLS5ClzIeHMMWBG
lbb8msj7xNYuIUx/kLFjXIB49mzIWK9dhn5BQM4of33jnXbff1edCjp+qo9xTHQC5fLZ+aab0lsq
L1IeAnfbpdAlSPdq/vngrrj0EYfaUfwMH/fB9tyUUTWwShT9TOffF1R4vZLU1XYMbL8wL1acpqnl
Q0pjnE8=
`protect end_protected
