package d5m_camera_agent_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "../defin_lib.svh"
  `include "transaction/d5m_camera_transaction.svh"
  `include "sequence/d5m_camera_sequence.svh"
  `include "configuration/d5m_camera_config.svh"
  `include "driver/d5m_camera_driver.svh"
  `include "monitor/d5m_camera_monitor.svh"
  `include "coverage/d5m_camera_coverage.svh"
  `include "d5m_camera_agent.svh"
endpackage:d5m_camera_agent_pkg