`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
oYtWtk+XpACzOXZ0QJ+lGsvU/zma6LqtAj6Pa5RAWJ3PMsEjNSyiPca/V915zehi23jb0ns96pMz
pMwSy/IfVQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PlChqoNz48D+PWpnD/OgmZZIdomcLWgGP5EYkzZPUrGLR22Mnh490obHrha4f/n97lwQlbGomLHh
CNJFYPxa/u1BCOLnggcPy3V2UqknO0lFeJ7voFJCCMw0DgZbLXUVGdKfLIgCLjJ5KJnBpuBa/Rgv
tyfS/+T0HiygsGHBGeM=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eAcsax5Wysm6gJQ0MR+ktcuTWsxU9c663x2WR5x0N8o8RvRpIZFZOpjcsQ9D5bXXYtRA2/RCKBKx
0/930f5eLZENSh04hwRys1qpwhLBf63iNgpxrdrub0YcEkxpbf2Sd2ra70jckFXTRSLmPrMGYkRQ
BEFNXYKwGe0U9yk6ZJc=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BZZcWESH2K1/ggFaZUilcpoq4DtJCvsVW7XhfjAIrgLKk4zl8PasVbCzlcOutpetxCGHa1C0O8Yg
vE6+hHS3wZWaTyVM4sAPUqjpwIBKgjDQadwgQxj2Iktd9pgIPGUErec/jPoLNCJ7fwubh1VIsWF8
rS0vN5oEDb+ns/BQQiI2ExBH8QWI+LuCpIzmg3kEoGszhQ8mGdWJ9NhyFn/tM7R0+9219oVwTNlq
QtXuedCk4so5eLKFF2SlXmQNMKzjntRRAlWaYjnLOmxaj1OHv1ElxdMR0leCMs8bBWrMN95MsVq7
KnypH9qYIWFsw7gdRKjRs5wILLA157BOml51Dg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eNcryJPUO1mr70/JQHnnsi+NQ32mN/D3Qh1OJmmHXPZ0h9aUBRzXNhndNaW++/n6bfpNvk0GhmAr
7CH7GSVJKSOVAM9GMrmTSW4L8RzY3+UVgrG2fKFmfmZVE7aCWmbOn737sVGDcLjuI2Tl/ArmMaVy
1Xan0feVUV/Dmutgh69sSjICauWl367osEVPtqYNLMgVn3gpHZZZqeM/L1EQYj39wbt0ZrZzEHo6
TYclPFGmxadXS3rPzvzV5T/sEY4SfLXiYwIV9XdmYqPXWZUFUsF74Ae9RCGcuVi4lXnoaA5e5T+v
Cl8UXKk2t+58Pn8g8Y/5nMAq+pHctnkBxGYjJQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GXalEFNXX2G1w7538XAcpC0ka7EpnD3rvZUfvaaGn77a2sBGvkm+tPWolNHUujJL2uOwrLHjfYvC
uOmqjDN8ONMI/+XEF9hn5uW4idFsohgp9nd2Nun1MktsJp30pldOwB4R4FhhjqQzJ4DnTzPrQO57
IT8SFQmZWru0kB4p/L58wgsFvLKsG1um80jI7JZpnG6pZGhQ6gt/Wx9kOpUVan4ypoZMT5XO2U9E
AWjUzEWlxhqqJYOTkaxSWJV6Nm1C4AiRlUU+W8KHKNvXfLwHYWdMWuB4EO6q7iXUCaQy5hbKoBk5
SFzOVo2wfGdGxw5zE7TTw6zULEUPobupL1pq5g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 565792)
`protect data_block
igSKm9nhVh1d2Zm6gl7X7trIE2mHxK+Q+Rjn+yUCPbY3xCJnj0ddcgPJNeXMatn7IlVXC+amtC4z
M/+0J+P3f8xJ8Yzb4VwyTmqiadzdDSGfZ8zWdsPqTOTPUIHAKbZeCcdlI/1f869G4CoDBvx1GaV7
d/4qNv6MWGsv1r7we8GstcKeu+Y/B1XY9jeoRmYPvqNed6HC7qRPpxFqlyl7UPZKLOoxuPI4DXb6
OO8lgYwzSuqQo6rrnVZKPfDED2tNYSoMX3VqxPDiI2flPUmS/njOIOp0MWQUI7c9Eqtsd+9A30wM
eQjt7dr3TwpUUFYU9WDdJo5hMRREQ+tHSgX4GMX//GfnXitFL6WpEOvrUgk0wMvr1vfh1YdCV0FK
PiqpR48k6xyZa6zrZEwHgoOBsWwmlfCST98mRHW3flq+SxWd2/8xFdKPSxHfG2o12Pyb1XgYxNGC
NrF6fu71ToBi6jGvKXoQZTaaT6TUy6HMdXSu8fH/4T2SjOyBaUibMHeiXf7UtmVA+2Zka13wbzH0
/fwSJPASvx6tl5W0U9QTh//p6OFkIs+keXQRChZLZYtBoEFs9NEeIG1RGEZQeuOrbpo1uIERjll+
if+b1wpxdeddnGQstqErR3fMPPeStaVO7fUWuOVpEEpVZY/Mq3VYTZ64NnUxtzmlb76801jvtYhw
PJIbuMwE1UDhqy5Hb4hovfLHhEoCC5+OKciR/fclNgWDFuQdEzbP0TfbrKGDBURFnY1M3m/R52cv
iK+l1QatZclnzfesk1oCVbQufyOY3lWBr8ujjLNFhnwrQyWYYO2kSttLiXrPHVuL4KTWN37E0eet
Z/FMtxI/jeNtBXzUi7Xx5/q7B41QWVqwkYpA9S6wcexAOX+b+sDsorouruLjMttqYedP2O7n3/4L
7VMdXi0K/wmMCoWfQyJhw3vi+UgYdJ2bBHwzECM6+ScrOzSA12+pqtpqdujyBUkUWXEoCF+c2Bsa
MRakkVqk+7N6ca1k9enJCYLjo/H7VBgUO1t6zGentjpvuF80ft4vTJvGgz9BtEyZ3UXz8UD8/aXq
4DCiq9Llj9y7U5HW6SZpdE2nqAPRWjyPCjWilJwespoE7/9qcHiXCwFesxOWiZDqMUTY/TReC8T1
RONOKMZsZyP4WVqqzU0Q8foOCuDBSqufw0EB2qpXoH+4+WXNQaHtEKFIMJrpa5+1RgJgC7YFU7c/
DdgnL84ixXLXHo85nqxDxEh9sF+4qLmOVJ0uRHIVy4Y3vJ4JI0sViuqjwLOFs9ylK1dpunPnuEQT
yBr5d20BvLS34jQbaIxpM2MmMwMLfNs62qNkdCCqHGaJkGQdcm9e8e0fSyo255XtPLAjwKWrCMOh
9fTGlxq6K/k/yBDSYjc5b72REl194/J5wt15yNa6HWBaGRAzH446kgQYrGflLcAfpRdgsWhofaEL
pRKeOmhzkGnUkZZHm9szeTd4G1LbCQLdWt8/zPMx2XtyZ4vTOw3UnSISYpca4Xr8KhnGDnzUhOBV
S8+7g4xQaQmyswmpoO65/0iUE6eHsanJFyxbolZV6zSPgLfM9s4Im1hYxJKlRIZrNa8Fb6vCXiZL
MxoqYczy4YHcgLbebUTwpyLLKoosLr7uj1v/WIpYm/wEAo0nzRLU2OeyzI+zHphbV+Yy3a8ziH7i
7uqwQBVERrMl7jdGUieaH0HqfLYgLAr/anjrqLcJu8rf4q7Sw8bh0AvDHKwT4AoeBud84d2QW0yS
+kItSd1dJ8r3HA3oxx6PiaN24v9x8oJ1xfYiXz5n9uydR+rNTdw8hrlnTegmm0bAVaY3XwQg28fx
xYZN1rQucPUGB+hAmt8Ptkacy5uQ3aul/MMhN2EjVk8iZCtbVfCmkaDTo3Oo/C9ewovCadTX1T2j
BRb0bfyaighlOS7bPulnBS6CpEgpg1e7YUmzlaVfyiYWgGKQemz7SHPkh7blHZG1P2iDfphCwqY0
gxsx5o5FojGjiZDi+O6NZ3V4fd0Cx9847F3LUMn9AXQ0itO5s2fPbUQIuK15h/dw+N1hERjZD03j
yTegajEF9aqTgVvvT65ZYbUc54esfje6BkxlJ0aLFLaYFvV4Xxx0knQ5urUmbLTK5cCVamienATB
+Bn6BikeKjZgjTYl7IJCNxNWNcGliYq+UNN06lETbzQiRDeQ6vhzl+GGksiH2lu3J2dGhamfUSru
ZoGePCAD1XXkhsE42OBtFZ2ISPQk79eNLt1o7cHoA0WFWTeFOPFftV576ziVVIhB6N9GakW0ufhX
fEyIXQ7vZ1bTqmausGyvWhf+LjFxiLYb8tt/rWDq8vSwWYtCjpZw52s2P3sbH3k0OMJitGf5B2VI
QCW/1mu07qyNP8JYXXY06GEDjaA0+aKVgUmdzfgbGw/yXiZo8R1fnahjccQ3En/ceCQuaVbX1VKo
tBUK0HkMlFKIZAiQ3P968bsM52RxWJFFKbciMzqL27XrYe3JfT6ExxtboSGXAQ/yhKTIkNTUtFed
rADzuTJliWPo8v+LloqnduerhOSNofifVEXcw16lDn1yPH60/yC1vXYMu7H9HJ1dbdrqf49T366J
Co2HCNQ3IMFBf24DQwUM9T5JNgzkDWLKG5+1sQBvG+vSOvMgWdi788eja9cUvAWZ8kjkvTKCemIs
IUa3XIE8BCkx2P4zDhVgJdMdh6A/hHTeaIFb74GGwgm4GAKRYxBu8lnKABb/IvoGgU0NXbst2D1c
5QzKJGr4PWzusOnAoQGdxMSi91jqDDV3XwHPlm+w+FQY+2oBudcLcMRQNPdx1bsi9HLDUZZxe94c
b0lO/Jet99f8OoNDXASTj/rW0e8156YF7iopmKntzC7beZH9tvfWAjoR8/CZ4HFIWw+bRRM1FtMX
GbU8TWP7XdsurF/3TgZi1zMVMZ75RUWIfy8A53XVicFA+suGB9ysVIlc6TalW1xtkiYX/BymZx8g
JIf7zb9QiTg1g37kyTkTsaIC0JLndjJmze5qpPeewtwBFl0yUwFalzbsKpWIEgTUUzDFRFw24zwA
sBAkEcy/ppXASerEgD1z/O+2ogKH8AsMnhJWQwTDkl3eYw7CmDD1O3KLgy+hwkRb/mkNCdumN/Dd
Eb8vL0Fj04lnK0RTn5eszurwAfR/cyp2c92ijgeFWYSFYKuAoMioneeZ5cJX0j8kvDlZySHNgk4a
ic7APbHEdQ/3iQQaX80Gowle9xSddripsRvVx3FUT8CqeGF8D/Pw9xP8BoX0ZgHQrcJ/aaX81AH0
zJnB1iNw3QEY1limjzwoTxggRsRgc/eQI1x5+D5GMWfrE8DNrTE67csjgr/gOp0Bfi9ssrj6yghS
osOW1H6Tmmo/PaW4O7BLEUXOsAFq8+RcTwx4BXqZIAP7eK5l7Y1u+/nJJYvYpXlp8u/RvQA6eoov
GYTni8r/x3g9PWv2qMIdhoKGoQng4ld0K+Q2/MEac8QkUEkFKC5H9gAW13iR3wAp19Z2FluJKjem
vpzBI/t9g8E3lR6gASs2nSkakZjKyyeBJGE078xaC6GddteBKNkO0pPe2T9gm4iq0u1KOlWWCqcB
OIdTXasC38bsrw1RagED3mV3+70YJYB5VZXWGyy/pB8t21NjO9e8mG6YFrGW2EVnV3cEI93cREiE
9jJThpyO35rqQ+vwi5ncW5a5xPNpDGyL4hkmLVYG9UrDjyB/PB3x58VAJpebtAv+mqYEwkQmfcsa
uIwiNFRYYJlecbYiTeutLkqgzVjYnLCtUyYyVii3efQpjrVybk0tgmxds4AsGeSJ7TGTIaBFS+CU
RC5xPn24jvMH5wu6J0AbZutdhVl6ylwT7EpSWSUAV+QmCQvp2QvLvAFSwFxEdOU1P3zGFfF6yBBb
JhnXgkKMEAfk6ntXAWNzFNPbQloMiYra7MDviUb7d3p6aNOswLixk3qyBUixLhD/Z87KCpl/k1zO
vyBndeG7gGxpNdPRK34iGkgiuwboA3Ot23HmupHM/yhGcJXtk8nsL1xtOFyI8Y5UuWrlLVYoJtn8
239d/92qa6fd8MWs5hq4nF6VUVV9M4oCpGOhpPIteo35w3P8lEbCDSzNBzjd5JDmUowyO2VJox5Z
54dxzNQ6jNcPHetQzf3r9agTBrT8+VN5pngFig1qRGF/jF/iizuSxRIyabJ9uEAaI59gPuPhaGu8
kbXNOnqOhKFHfCOWfZtmp/NNhnAQ53SrsVlMV6grZltdDwMl/+Vnsq0OzdcrqlbNxq0ZOkZnqwG1
JM6MpuwBw27RRci4N+75mphhWsMfpYp+GDRdO3UwjB6/AtTao7FqsEL96vkFXS462tngnYJiacm/
2J+jkXhI0mE+j1FWmByif1/UtFEFBWZEQJsCU5k8z4H09MoxaGawVkREGyCpViiaRC+EzR8ucfJw
NqfhNHIUfD38eBmzQOSZOdjnoNYLsctnf8GbFgVxgnAsQpuBn6IY1CGWN3hI2X0xKIJYCAqcY/w6
3UYNIkr69WctOmOpxemQnna9qde/B3HdU9vFbCKR6sSY+UWVZuZR41YVMMz+V19oFScR0SNCNCMC
vbAaMk/L2guCwTcLUCVQcYT4q262t0ztEGWemQZsgTcpI9rpoAt645xOI2iR6QRMqefubYCwLbsZ
2pw7d/MTbni9Ife9N74mu+4AOJQeaFPxQ87q68ecLsfeTu0at8G8OATHG0PPufEdLSmDWB/Od7IY
gqbwQWQwKHxRIgoAhJKrweBHdxjOmRwnWFOU7ORFMpLkeSvcTYQ98tHLrZbDLblLquj+RJrY/xgD
cV955xl4WDsmVr+MbMGdUlfTSSkCr1xcwlNcslKMXltTzSoFcStAUjRs4Sjgy28rs2cHVvKfaf/V
kER9xmLPyV8nMVgDUrzoVd8IIGu9ZM+iHFr/Ndbg+kcpP+rzRzwvYlFmXTxz8jXedHWKS/QAn11S
yIlD2mzX1p2svytFQzDPjPZXNVDipGLaJUIQUU1pFZ9+H9nuDiKcPl8SUfF6YfY2OcOtvpKCKHhf
UCIE6Mr7SOiBiopagRzSPB6GT0jHoyxAcgXuBpoSvZKFmTSEEkMORTRC1GDnKHhlwzp6pc6HxMRG
vNQI30deis0zlZJlGfj8NqykS+WjAcf9LjLYTJvo7GDRCjJALdy28nIAi/EohkA4eVAb6wvPxbwc
ZG2Ng1u11CVl3s2/XCyOjMDT9ce9Pm19udhsVBKP68AoSjq6fb0CSDvAM/qHjRKnJLiCC2cXVMbb
gVQ7GuUtLAq6WsUYK/OyYF4RGmaTAIoUfZKeYxJ1EvAynYVVdbtjvJF37ANLwrFkqI3rDWs/Al0c
mT64+yru56nc/cbb1mffF0eiHiVPr4qFuN0kL49xotS5i/LqibE9grTGijBbTgnRXWp/m2l9UsLj
I1/aui5L2Qp4Y1lBC9Dc6wCYESGtV8NZb5+F9CCS/zdW/Nf/PhU0iEIZe6mzZejZ7yvh2cyg6pLq
Ggq9DVhD0iJxL1jlE7kF6AXvIeTZ0Saf4ZhTLpBoh5v70mmwlT4rrNNFXB0E05nrnOpmbm22ZUxt
XKhHZry4UJhIPppFwpmgCi8aXsOdvGM1fgJ8ARtITycPWh7bmOH1wZ33Hn73JLA3ZPOqAoOtpP+m
F+3GZy35VroeiPRUNlhhc316xNbCeuCYJuF3xMZfsb+rY8hCoJM6bOlXL8xwzPZuIyqRi4kKI5Hw
QFXA9QTgvhnQ+RcufpCzs21TThBSIA2DG36IPoJb9mKulTza9+HRs9dIkbbe6qN3d0jMzUCoDrTa
u7R3sIA+FHb26AqwqrXbwI83y6f4476NLp3mqGuTBsesGlZO7Bq5WWUfNJfqvRfz7ZkcrWrJYpAA
RJOQBxU8AsOtPGF5UJrd4OhuEFfitQa5CQOrMFd6yurrTR5Z3qTrTCXUAMdM+Chu/ycVSVjeW/QR
Aa6CcuhJeskdAUVU05iUupn/blVgVeZQjAqAnTYRAWi4rxkGbzDWx4MrV0y+XvlSlaZK/a7X7Tnn
oiBIWs45JJ6LIf7Hk44Earp9mmMUV0mUwKRf4idiR1kg6771OSBhJ1dwivwgxsDTaejzqOH1mEbM
fPGzS4NmIM7gl3EqZUQGT6OjwQtf4YmaegcYLrEyrRTonQXWHYNAsjDCWeGP4pRi3De38yBzq3Tj
yDQZaWt1KeXg/HGgj0jhoTjNGbNmoAM9oA0IPg/+iKWiTkOQydEDTI/0Pl90YKCTfYVoVG+XarHZ
RVyfB+Y3wUNMcD7yVEmtMaHNbUxXnVTCx29eiW2yjftY50FIxO8W6GzuDtADHitWqfUlPCTjire4
M5k6A5trYQkUInrGsI+5L02/JXdKE4WZNqZnci0wy/BJ74zlS9AO22saSN6uLGYe2j+FAYQ95wNu
LX/wYmatjDwEnrwdEVNuxXMvyBa/sKy3lg02g5iVuSoVA86lgpa4GWBf7Xge41gJgFWGNInrYG+N
BUIGNTM6nSKTc3zAhXD75g4s2wK7F9Cg384cXvUoa89Jg4CoE13ujU+K1ItFVBSgfB4zy61In+pk
gWJCBoHpj/3F5VXVGXouBJVhls4YIaqUZjX5IrS1r7dGgEiTkjf1eBzQz0th7CuOSvEH0EhpnILe
KxsYzwL7niAN00OBQbl+hzjT7Zv2/g293KCUzKt+cTz4p0FQmuq0FuTImekXX2q1OT7WFdXj7Xf2
2zX1PPt0CtOTYOLrTl/1vqBLXNyH3a2qtl3UxbZlLWbsamtu6l0nUBauucUflgknQARPvookAPbk
AfZECIjs18A9eIhxNE36Jbct65RzAoiOLxbh4SJecsyfx11uQG4CufiuXwAtrzrXGGm4KH7fHtCf
0X6pVPopfxcFum7UO2z52m/RjKpsLJ0+nrRL4kjDbKzSiZ0LyDBzrI9v/6QZO2JCyB4kxCGfce9D
JX/qyXYNMXvNU15f+m542kVl19j6SswsJADYJkGcjs9vuzQuxjkIsO3heM6FApG5YkSrBT9rJXlH
uLKGrST/FWFZ6t/d1XxJolDlL9kXt/d7Q3mNwBnkZ5dTVJ0uExs0JOvimaav5IKvIiEOtoSSfV4n
aR6jMizgkHJj2N3k6DgmQOx1NBRP5sGNx9rLpqe4m5Z2kRVkPH8859Ge2Zlod17Uq20NeVE5EtWg
vSFScSs7pOfQ2LaCHWQxnnsz6ltLVoIJxd1rAe0tuF2xqUi9ihLYRvyejfYDIinOdSujw8qzQauG
LMi2/8zeFYMteIogc9TGIif54CBrEIg/PsK6hH7XCORwrVxb2MKY2JYFmw0PTppw/LVCvqP/zDPf
XYVfy4PjT4CKOcxtTP1VLnEgIeLs7luwd5OEm+Q1MLmQp4Wa3WRsU7anwHj+vXXDbj6coScnwB64
TdbnONFZXilbmJ4BoEh8XwbJGFPTSBuWrMxwB/gbuKRLNKPS24P3zDgyl8DlC4umFp3dKkjKWUBZ
iqn/leJrb+7YKkX32oTQrICwIp/Hu8lUXiZ/ikRiV8VgfH1J8Z6VVmevliyY+S/JxkHcBTqWVaoB
aTWIcEMdaLQlZqzyESf1W9Ci71TPQUJ83TmnW3dJ+0jXd8K8jvq0IiO0TB5PaejUbdyLEqYRL7Jv
ED4XePoIPpqSe4ywxbLHCPP3+2iby6ECjp24ABkv8jh8j8xb/ZeTFtK0aKhTAOJuMLZlW9hMIoI2
naP9ErAKZLeBwtl0JDCqS4uIikxTsSGfwq4RaEfkp/c/99Y5HLrQpXTVwWogdUlD0boV0W6xGqd/
BuW0ch881d6MwZIfuYSUYwduiD2NpoD5MYIrAKZhatLCo4BrMWozTo2cliZK9bXS139rMl33GoLb
jJSxa4fx3YpdgteqFIeAxG6RUYqiEl38W+0FRJqY4t+gYXd7ehDbFesfnlAiKB4IQ9vJDgThHpPy
9C5wsBAayULfLFVRX9jjJHziRs4zHJGAbFcDC3NznIVlH0iXbnhJoILpob+c8qzIcHQvwYUtAkBe
52jRl7usts8IA4mPuSXvfsewpLppzh/z+/hPyBtc6emRB5gyphdC+0lfwTT6JghMBXBGbzuYdzTI
o3GNnlB60VDYJraDV9EBsI88mjOMDRKZIDJ+VgJ/HW7TJuiEKMpwTPDflTzJqlR+gTNJFXVs50Vr
UCddwu2eTMTbgpFEp/+lrhMkyCD4Y07FSk6ZPskkzmkbG1P5O/z4ZyDPT5mm8W+Dj/9s5QBiSm3K
w9z2em31xjdBUtGLx2R9Bav2k8oNMJPNlWnTk/TtqDwBNE28cUP+Vpyuv4+D/ME/1dmlLIWN7d3I
puoKDvVe6qGCzfHVBW7JG/E4l4nwmpTL9zu4kPMj2lCRQO//XacDROr5B1db/HRRe1fO00xm7vDy
gizqOyCH0f79ScTwutOtpnqJ+mQ+FtQprP7Bw6xAT+IFQM2ZK0gwRcJ+FhT2h18dO9g2Nda+0t7A
GuAGisMi+yEZjeljilu3Bqe+cufOYMiC0Be2MJ0XJkGMVCu9PtpcKMFXe7XVuOOyYs5Z0GviK/XL
6RszvI3v0un/r6nQNR/dQRBZdBnnu8eaYcLlmGxYkwDrd8LzyFt/3ItuIQthfOB8Mv0QEkTYIfW2
T6WqybOBXCeHZtDyXJSQMXr3GCqHIjxjYv639KL1gtnYHS4aJiPHKz/I789wUHurbqMFpB+Ey0Zl
a2yUjvNi8x3RSdn6CwVFYzCnLl35LYJ+4xn7KDos+5bYJYA0lK3QrB/KSgyp5lTZbcKvhck0PIAH
BhERX96NhlBEYVN72ELAi7clH4pvv/S56BcPHtq9AuTErctlWTgfPll0lTic55cLfPirv6Z1dA2l
sKY/U8VqY+59M1DorhJIzVuxQ4giO9O9PJIQftf4m/PGxpcGhed+kPVjzvBAEcYhC0qxfeloRCQL
JAmNU0NN/U9J7D5mRhAleCe++L7TM8XzIDJR56DmI/GzQoYEUd+f2SA1VioRUpfKqSu6/osiOZ6W
J29HDc7WhE0zN96q8VgQsLSYLVmOEkOn2TvleUlrhewP13wR+EzMw4ODtAxmJzA/2WSuXuMBlubs
Z4c0wZIlKK3zremQmE+ZWsn5yFc3L98vcM7U6N53JIGsRvnCJPkhMV6gZfUon7hlB+R2iAuy7n4M
DWH3n7QjLVCdJPfhfHpII6FjFOUB1BYRUYZKEXWjYiXiEzFaYqGf5bv7YRC3UkKE03DwMUowQe/S
r4RnC+vYbKg6ODofpok7E+Jx2pVK3aMZzWgJ3PVefXcycqhueu88NEiHl6psYEbYOO+Xk2XUQPhK
fTO28SFrrAefJKydM9nLdBwosd7aAvrbRGBwSHV2nN58FvXVnOWT0YVzMC78m4i3CeP1o00AHmwY
6Lqq9Xx/dT/WbsD4eNqSN5UHgLzpmwoRZGbTQOOpc6gQj4Hnoj+ApfIxjoh+yg1n+M9QmvjRRQ5q
thYQb/fkcnwNsyINLshTNq2PimLMBSB0cxD7c8G6Mow4cGm+kacDUAnJvGBFs59Wc/Gh7Gz+o4dk
T/0b3qMDqyc6nPq81JABOF54BHlMmt1HU4FZP21XrCo2HYWTiYawHDJNOjDrJLycJ6QY6NBOTpZm
+opichgJaqndPSFvv77AkSrIdvdIh1hcKopZksTASYV1irxIk1OGZ+ATvqN5NOZc4KxpJ/H4j3Yt
zdQ9OZg027RTvDeKFVGFQ7xo9/1AsCom3caTGgZ24aB4Gm9XdRCVMtlkZCYwygDQynn4PiUiHXGR
gZA5tY+K6Pwm/mZux78w9fKaJ+9IFkuHCpTJFDahj/Jxquc5qPJ80XYjMa6w79EAkH/ljveJydH6
DFWPROrfH/nVVZqQQo0gdxBeApplPrkYAjLSlHGISlh/oasB4wvb/F64/s4LbbOU6PPfYopRUG/o
tZGI/Kv9caMFC4EPBg0YBX7Ilk3zhm8hMYUMuxCKZlK+X3E2Lv/R45OHBDyz6CzjedpOmf3pLVGC
1N55Jo2ggLDklz+KDBhL0YpONYe6a8DfuypNTChgX6VV0/IcNDz+jObU6q3yvK29cjk4FL+WGaZ/
UkQTl8FVEbOghV+rK0Rc5Lh1H0LHBMIojTP7NnyRwl2+4YCrZAkgBfMyEPF997ZO6Rt+Eihy05BV
VuKXMktjjD2fJDxFYiBizwR0v4LKeF0N7DgBImIE7f2Fy1BnglN1yc1VRe0WP4T+1JtW9tgSxNpK
m9IY7aFBfZNnORWu8otU5KkcJkW97E615R2VaXKFpAM09a5+We7G8iTL9NQm6/O9qD1RIpaI/tvF
+UmpYaNLE1BBle81W2hWG/d7HzDSFRK1TbClQM5Gbu4s+Xy4jE67UHzyTTzK6PDF+2cdnd+WdMtN
GeqMoO96BjtaqoyCNt4HuOsvhLWQ0YFy4EQqsCEKwAfwJeICSkcDc0KDJuJYipBU8rcUN0aA7U1/
rV4snCQh6OWyvbp9nXzw4AHYOFuUIDY/w09ZfPl6Yk/aGsp1W0pcyDm2cEN7Pb47v8vy7vm9I6FN
BiNdupsZNMEl7oA0F9ZaJwjuVM2lupzWBBy6rEBXKvTDcNM9AwVKeGZDxjTEQDp1OtvriqHQGjf8
ZKUtU7vL7OwS0iWxPGPMTq+ReX2m2zckxykA1nVTZUoiCq8Eso6np5RNzlNHjV6oepXUfUtR1d6D
YKUKqlA973wg0A5+wCHhiCBOkKqygqZOhvi2Lh6/BfN2cfZu2Z2BTItTQ0oGj/ozCGU62FWw+xY/
OyKs+LOHOAZYk4a46GsxGBnBUoJCQ0tqNlisbCWXnsHgeFEF+58TfMU8VrB7xJ8E4TITTVGGAYOQ
DzVGbLgYwejlU04I0lB1suo5Nm/tunyP+bPR17NporZBXWJaaya5nmWOxhzKZV8wJj66UB68o9NY
BbzSwme5f7bJ2jdg/zXdoKgsRdCXv7AxSj5zjvxmmPeEuETnTezd7bnj+nGLYt++6tl/mmnE/HbM
CPQ8OKKdduSRWLlANJDeB2sl34qRosg+nkGy2vA3bfsDjDMlVJ1JytbNOjhpoFX8ivKr2jpZhdM7
K1Knpznf7xEf+wxCFWRdJ3krzhQv9e0SOy14EpLRApDzUUZnWFnPLeYoeff+sorZfZLSu6GR1Imr
oBfeCECLCAhL0rBzTM/glKivow5pp/peoNwt5z5i56/BMqJmuoobynLe7QXJOqOBr+s14MSCggul
Q3E41B6ms+0IY/Af6Ir8WXk07UeMSQyQfo5PCmjelgVY2kg4JF+RDiGLdrSD7UsoEHxBHFvbiea9
EuMZMXO6/66CQTZN2n7N1QlIyRQS5uoN6MfgYFkIKrI7YvI2PZq/Kjoa+exuoIjK3LMCbWRslB3b
1GDSWplXwC8a74kj0z8PJ6kOyoYIgqV9pguf6E5HwMZT6zx1O1gd+wfQv7nhfefXRFUCiDCfSRcZ
veOZxt1pWPHcMjmANuPkh6XCXTF7WFFRD0Qo1SNl3AuKsthTaHcjZbNT2aGTMdDzNQ1QeE7qxUon
hkmVrWqa8lDzvB6/qcQwnQQGI7jl4dNvxn+YCMkkUeqNEFjx5zviJK/jDnVurm3Npp3DrySKph/a
lo5SD80VnBR989JaTIeaDI0v4An4Riqc8gqMpJ6KiXcyYQnQRDQDz6F3vFC/qKC0SXfxpyTYzbaD
NZClCBCE0cOit6lJHRM60EoOI7/ruZJhDi16i0DN6D7TDrWF7HCPSEehq8+FAl7zO8pCqB/TZkIm
8yDQI3Zp64EZvXKRcNFLUJutvTJn9iBvjmvyd53Ignbo4FVrFaiCCpYJpFQunYZKHCtPMR+ZIr/E
k1xupBwjtYW4MFBhuXM1ILW2wNSIdC7iwA2rBXW1tveXtgDYvQ/Uor61RdlAX17FZerL4NmilnLj
CeSKkH1qi4jfhvb7UlK4cE+9p9BgZcbTBQB/JQ8/TE7ADFF8rNWULT9DSnqPEWoREgTdyDR+nwxe
3mKpwENRgxGC/FzPk7Xbl0ypgjTqebDQmPoJihXq73mkSIzv74zDgwXjx5qvwIiRjxT1VsDB1IVS
3iJ6tWVnbUV5/Kvoqzy52jmgzXXP1Szj0ppLAK2i8k8oxpA0N2b0f9wKfqCENmR5vvovUQ9XPnrP
DntRY+hAD/5cdxflIpTEJ79BLeH8aJQugkhYuSuZP9pfyUywtcaU5syqyzg9zCTWTUOEAt5JSjba
Rdry3FszLQ8RnPQWpQSPv21XQFCEfHNRQBSu0qEvcbYH2ox4Xg7CnkswUfv2R95m8LrDktf150U6
u/UVLXBZ0WX+68SZepkR3qe0egjUHemOM4g1zZfQWZweEptmiZwNxu9NN0lFP2PhgXsDy6HyK9GX
KL6CedAn/fnGDKIBhTNC6YFqWuJcijQ+mywQMLnqjOXoU6jbTZ4G2u6cbDvDdhUnscbJa22Js79c
71oygsi41wgm4TJSbqTXVIHUzergBQv77j+gfv45VjSeB136Sj+MlAl1QPXRy7PEcZPteUscQDPF
Aurlkhv0cQt8r4NejI6vcFdQxv3c4thkF9+GvGhGd75aMhUI+gnQmTFMws7Cw4BIUt8DErflM7nJ
sZ7QSQzyvkBO6PaBRbnfPIyE47gnJVYHYhRwRQnHGz0bVbl3KchIUJn6oB/W+4xJrz+M3r/SLy+A
7tv3eUY+w+TkQVJSsP5hcjKFSuixfBRAKMwuNulj9QM6BY08CBZPcTYwJdsr2rhXRkLCSdDhLzwV
nNmG7Wnz+dvEvtZDcF/OUkWstTjeTyoD85dnX5BvW/G8JMvNU2P+2yRVf/RzVUadkY04tIlzk4mI
Fw5n3jQiKMmUIPkcPwXrsvpcRdtk7NnYYfmqMef4maxMdTfUrHomsOU3DWlQz/+5kslJ+g+eY06+
xoHOPGUYsqWm4P9Rf0Nlj8zUBXto1OLCqZXdfi0DSNdgVYfdwx9XbnrQlNe29r9KqHhxYDRsqcBp
tNwx1OnKB9Vj2Ez/SxB/VMIrMtiRBBnD+p6cmjsgE8QhYP/pkqCnU8dk6CwVC7ccK3xQhdgCoRD7
kxuHphvjpfzA/hmHSt3bkq6EkF/Tvpe3On3PJqGwNIBjLK2l5eDKuVRC4zAe3FvwHRlFAJjCym4w
yiOQ/4rjKoycDN24rXYsKxnJEW65ScgBB2orvIxHgS5H6+5fnXVrtQ4MPCow8o1dLH9gf81cBOLy
s7nLxGXqDVD9dsLH5VW9UpBW+5CdH6d/8wiPs1MA6WTptK3JHwRXSP5XEXNLofnlReOZBKDBdlg7
FYcQ8iUUr5DjHYq3P97jv5D7qsHXdRp5W4Rygox6yfakLFPnShis0xTPBsvdjDmjQ8iVmLNTchE6
AQQ1EArM8db2m8uIPSNbrT9CKJH/hnGzsGox2n/lry7yvp0K2QVsssvrF+t3BQqOxvWke2wsw/lr
ZSTNLwk88NUr9jFKhY5ZNo18GIbcelyPaNX+9hHTVEAgeXrbQTBvBZ9JplVd3uS7mJkgYoxUYnHd
ex8z84BGGMa0j57CUTBqR6NfdvXwgM0x/BmwpO0XqYHEPGjNQtyQh0NXt79+NwpSlPMXsMiTEm+5
oMm7LEJTUVskQDtYMPP4y22UPZ0CBb6q2gEP4lSjpROoR3tosrB8e3tUbz+XXg1FBMAV/LAgWhua
SHoZ/yW0HYeCPKddQ3b9m4ujeJ+tp7MVnlxqTEfRuFkKJ/9jVgE0AItXbsCSsvKteJPDUhqmMnpp
eV2TY7AegJR8rVYibqNo78y65FUeBsjto0wq2fbfu6iNi3VY69NvELlr/Jap/tzyvnmLDHsRZnzb
MYFowb10gGNyKSMkpLLOemUj0Rxxj029plJHPEUiL0+A5pO4oJ4JOwAtM6donqq8OaI4mMSCBs06
pFpiUsfzqGZgCKMtjQCEz7dhmLj/Ir96rakf/piSOEoJwc1GxV29vFE54lTAr8nbWjmUymFAqkWS
7a46GkHqtyKS3vIDpNEofHDjGSrE2vbNcfXq41nR6qSd5G2rSmA1fvc4goacSElArWDMRkqpTdsJ
ad4yMVzVGjAn3586EhSTb+aleywhOS3uqYB4xsQ00sbQ2tvJABxYTCnodXODkQKH9D+S55265XUg
FTya4dIYXXCtrC5WQO9rTMajFi/lsBEYAgx5Hgn1E/ev3s1HyQhiW646zGPmXA+ICYAKTd11UPfM
i65ZyPBbL45NnEJRYj/lmQoQO/bMdFHZHst5wv+yxsMAOlNwbKzxABm8tomuffCtexM3qcOmEFmt
MEUa3QiAerJzHIpIvlGw/TkXsfiXKDKZvoLyidiNxApdLVlGb7TjUCTtcVxevGQM2aZOZxNXonPe
CkmTFh9dFFN7pnbYIU2jUELxRk5u/ekyzPzusxb+B0lWsxQIAYy+AgGX7z/Xo1sWTIi+Ikp6bxpy
/UVz/o68MG303S5WMvixc7geBAYF318RsnHF5BHY0I97eH8Mo2YH9QS+3V3arVpRy7rqJkYT34CN
075JirYfnlwZMB5Cf1YQt8wv63mDKtGzKU5UFbTnCeFEv1rxS2U2zCgcFxl4i7wpNeU0IheUbJ9v
thD+DqggGD3oXXc6FvBx//PrNncwDhH4nskGDqBd/IIl0B7zP2nD1QEsjLzaEqRCT3fgBOxJmnsz
plysJV3lwLChvktjwwG+9mimbZ2znABC/bLGonyoelRTGLUdUwxEMsU9GEF9XEYv9+QpFtC0VOwQ
2wbzURlP+oW2NIH/0fkis60DxR4agoL+1vA+id7BC/OwmmB0TVbCcI2MHuJFfg8mzVS1nZhvraHV
+jYfAjrENNzYbWP08PX44dg3DmxAQemr1wge6WtjKEljpSwbuQCwKYX0+U1uhRGR7TevUeYvg2tk
9mTzshQe8NYBC5NJC/fglqt/lZfThSUal2rE6r1NpF4UG9i94HFOqSNmCPhdmEa/HIb7VzSaI4kL
8sPFs+fc6xrmz8WxSFsbvrF4HbQASroXhRSvzADbk2PauJUQ/yevnUTgrLg0r4DagRokaulhNEVj
okFTXBAUVXfuxji811evms630UJBTdnXKkzhGqvmjx/cHAdU1EWjRJSBuzf1QHo9g2vdBM9Ramvz
0E0AuRO3beHNRC3Xaz8CRKMVA0pSxz9CAvriIgr1ZPZKjqVRJl9GwU+cg6s5lw+bE5YNPW4htkpX
SAfIemW44eBgQOw8QRCpRRI3u0faKlv9tR298E1VqMqeZuDTJf0R56FVAgQslsIBDU3m1uSrbLzd
KP+ADFxK5X2STkdZdkWBsGnYIEz1q/McArczd0lUfGU/lC4VV4jURKU06TLCZao4y5qOzcI5Z/sK
E++13V6M3BnPLM9GNWPQ4IGMDRr1L3yZhsXZsv2qr+gYpHCdD1J01gPhfm4thwWi5C0hgToOrB2F
k6QvntVoPjbc+o114bmpSMU6pahlfoYiIiSlK+c2uxSjZKFkQuwLw/7POMG5YOm75jp0laejO/rs
GeilysS4yySmqrU2rsARlUX63oAyjcv4R9lrYEAxC4jVfMFF8KJjQu0cVX7I/qextsr6C7RrGPgy
aiS4tqKWsYu1/M2MUHCPRQpkT6ZkSa5FcovzaWyrsYE9S9Iq2NJ4GnHUE1zpiUGtuDlXFbGQgDpM
urChqHcJXAABRs34EiQTmVwRk8MduMp2UXLevyizv4+S/8t9IbDNgNMzHJRXIOqwIl9p0ux26AVt
N0+URY721PdDdZaXwIcfXP2/jt1S2M0gfqUgBp/CU0Z4jPIPXOntFRxiKxLBBY+T5udyDvkGYJu8
8FLXslJm9u2EEF3+/CwRNMZbuhy3B3r/+n/SCiNwH7DtuGVDEbFDVqPuahDp/PHz91yQ16HkXcV3
LSKjvZB8amMNLPmeZAouyYkjjRy1MG9R80G7/sE90XWCosDjmwwQgGWPYYFmvTe3INPGdCjCFQ/I
g3FDkstNBOM++Eh2YboEh6DlYkSkxIwQpTVosbt3yHrDzxd1tVwpnJQ/NhpA+AxpdDIVA+VqdXdm
BNNKWkbWq9qsb7RyF6V32kE2h+Cw0nEhXWF1mvqe8odWeeiwUKChgnBdbNqYRgthLoc2Xu1bjYt/
dkvJBX4Ug3zuIM2ikMWwbiaLplQw77BJyTGsUIdXiUvQBITFyTt00PpsiHCtmvmdqQcTnfBssz1R
LlOOW5der/jxGWPPJ6Yl9Rp82LmlaccVhjxARxC2BO3w/fx3LpEPfpGlrAu/3O5tOPNwGI1RTemW
v2PD2GrJI+VLck7NLWPPKSm1xKkTtdKfKpB6EDSdjgbYQc7Vf1JTVkE2Y2yak34zdxTFTVC/ZvjT
RwLUylB7zKYV9oqGkAo1PkDF2JzbdJOk3NH8vjVr26bDg2CTWD0KT1hzedBz1bQq6VxpNK5zgI3L
efqoGazZ/nXoqsPZX7OAX+wg12HJA7WNupnS/RXL65EnN6B8EIFOKmysAiELisKTRJ9P8VU7VR/X
wlB/EP7tktkiygHOpRkuzUERCXMyPl8cLmVNCEyi+blfVfJgr2n7s536zFMJco7/q7z0oW4Qj9b/
rNlN6niv3DPt1TdUfBefEty+QvRjbyzFPdCJsKnWFP+sYYE/4fYF8QZCpgD7N50HNGvfUNZ6cVN8
hvShCsHhZ2XynyL0pfGXEaav8aZtkn713kFwDq0/VB96/ZQ1hYpH0DrnqKpMf+7RM6a8dpe/OimI
1Tq5d5na1NJaZflu/Lraya0B709KJE28Ukxf6shca2vEVN+HH7YEVFpZNwH3Lw9rn2TcGT7LTQas
q/pnXjQ3KXWg3iJL3EZv/99kXiQ78rFAgXv0CZOmBxQGK/A/TbUPJSgsDNNK+xym5ViKBL74O3Kv
0gmR2P3D1HTJF0dXXTG4mmJQFzxBDO35Hpe2+tLAhIRqkeFFcH3tJPohnGf2PT4it6tSvq0z8fbF
7aJHx8nAqSQ/cpUnOYIONJJmupijabOhHSvLoFkBLoKIN5xH/uQJKPC0Z5zqHcjfccVjcpNP9Tks
7QLPq2r8raa7ra/zBojy+uaXPytkO9en1GJKT7Ubimeaj4hYw1mt8IdFl6kIjWMvCLGPsfiH3uK2
vH+6e6QK0Q9qmhtHANXp95wD5bToHJQSNtruz5OPJoWOw9AhrBSQFs3A+Ot7Hzs7ayt3SG/x2ann
rGD+PBpYWpv3QsifSB5FIO2iZhS2+4dI95rEHp363RQiNeLXWcviQoy35hgXLl3A7oFAxGevRfcM
+h6ZVW3fY+lyQdZXTjxmphTS5nCKRCP/tIH2u4k2WoQqukbusMIhrMtx4QX0y6BC9kmUOSovEfDD
ZuXGGIXVJvwT0yvG3o3kU9aHlR5Bu+eRGo1QfG2ZmcFgoBBM7TXHKzR4W/Z+vuJD5N5aweR+xNRM
kGjPtzZWVtqYhG5XAkdvWeR9YfPPsEmNwAaF5NNBccp4Y5zoEdDIrg2DRMrR5y0GDoEvn7lVTb25
ldo+tHCetNpC4RB2MsaMcH9UdcvNZp33iVP2qm0ldu/rgub0wavTbeIAWkvfqyX8uqpJeAAl2KYa
5xFtjaXpfaPNsFiUOVT7ci4FN/951DqGoeTQCmy1wRupkAHMxyFziwsLYa32d08FQztjtzPdcotj
u7dOpvu0w2CpJto+JkflfPvKZLh6TcCIZooMkfp/N2f1gX6OuKGQHYU5QHQnBIlu0WQ8KKCjZ5yN
G1TLxeJMQ1Alz8qznM6qR/GRF/q4FGNOWlCqSqur4ds3zgOF/J4ix64jR4hvu1ZzRch+tNfcGyeE
fzi8E4c1xAJgQIzH9XQkDdQRj2DgdBsWDfIT9Fj6+5BIUqBPSGp8+QQ+3w/RlOylvcZsv6J4KWnj
e/+mhHu8+RKS1ecXnexMueYrnbNNOKfSxl+KwMv92u5/J4V8SQTN8fkpPiKF1+3xUoRpd4Sy63xO
3EQGlQH0Yr8Fw67sOzchuT7Yj2tHvguh/gUU5tEkZKSUfvifBhutZxOlW5iSfGJEFble2vnt8HS7
dPsq/x1cnGNCCnN+lMHSPvs9dp5FoA+rnWsVhSr7bFW7wVbPOT7FYg5luWlTXmLB75u/s25gIAuP
laYW8DMNnTrevCbzYaJhn0NIzHdDdGQSMBOwUhckOR6U/TF6Ehyb7aDbgDowCQAyG7downiVeG2l
JZoGQfWGdppB/4y/PwZKoFSEHUYSXnFfWlnY921ToTx8QgYgjdbMM0LxUvcYrcYps/kdeooDCMTF
ygjRH6D9Kj+aF5UcVv6+93v34LXGRcY1EE2lpGecWptTVrBguVY4rztwQAArnIZnuIH6EHc9cKYZ
J50cUtnJEpMK8TswKxqzNCin4MWE50TwBz6s1718w98y36NfFMvCIN+OekMUOG4gHEteU2Fs5fPK
sCufeFSmVEruZCroIobmc647MhvR6VHWPUJAcEJI3WeDZ64BIMP6hSdqrC1rbUR4N7CM6NSwDcmK
SWPy9jAAs924RtLD+WlMPK5u31l1+v5GlDXrJWaFJsDNc4tALbOmmmbEGVw6Q1nxyrSLFZmbjODy
J7Lz8C9xex7aKHWXVwwplPjvkVLP8FEhm1nSrt0cYyqqp5UDTUFGM2UIR4qH1LyRvlsGHBSIKED/
dHGsoW5hztrvSrYUuswMc89FowqDI6fry3itxrYlMK6/0/xzZFtc0/W/YL1iLAWmsU1o/SSsAykc
vkP7aTHBqS97+FkksomTshWXEVeZasPBIC171P6vcCzFtSyAss3fyhxZmN0UJVQR+H26zr+rG5GK
ILwrl0R1RChvHGDt+Dg2YIWaunDY+OZA6LNmbCPB6E3aoKGgZkr1fOmrqVMRpRAyON3cSw62XGmW
FrjjfctAMi3yrTM9LilS+Fein09tyx2sIUx5ln9WBdnoA7cDuehDMYbTD9wybJ4d56eMCBENwOak
Saz3SE8fdMByeFhaQr74YHTElm2gCIW72tqXccjVXyzbPBQ2sUYrhqGGBsBHfBjPCD9CBNVVO3Bv
H4W/ZmNm447KGT/37kYCocXG1uwxBOi9B/h/PbMu6BkptWiUPeszwi3O6er5bdxA+JMXoTFaJ3c8
StLeO5uSG2Ef4SJYzSZEPD91cxTv3oKHdSQSZo9HFPKcHywCSnBPSRBsBoBg28n0+rVX6583gNjB
9b04ZNWGaaznkI/gGwlweXxCvQ78waqZDunUKiqSqBHBBapxHN2yaxwOdCNvfD87GSkMmvHc+3BO
q1X5R6rNbFHWJxxFYEKQVrfsJ7YcUVA+3vWzdXV5oZLE8KyyHwxSe73s78jSQ4UmKIeB/dDOr3ee
bxSMFtPyd9tyT8RckZv7wwYT+LBxQnC4RV/b3hx2eNZ5PVzb37lwE9lY88PzIA1e61jvfr6ZqD58
m0LPi70QwWO6aEEgFRvQeOuO0BqRxJiXi3SOHk1aX453xhjoT6Nq33Dg95lJSufP6jhJSnlTRSc0
nQ4HsOTHOR+0LZuYexSH6iLbGbC60xcyx8qdMi8jNMbE2lxOVzypkOtKc6kAwwGenDFsBHHDW4wA
2nCQUP94Jv5lfOsbtNajfGkuUVQtjVil2dUwJX3Lizb4MyiElV4QpKQpyaILWIoI4ApWf9wmtz/y
ySxLJRza8243umToMe5Y+q0f80ST4X+X+cZ4tEa/uHJGxbQnK01PSNCI6kXcAlcS+xGQ7bhffLpj
zaK7hChME7Kfh+iFxRwwc01bcXklum6oV2ONTdzPlOLtl9UOm5rawhyBA1mDGTJnusHSr0DIxRuu
z+YUUrNNEcQ5UH9mSdH5iezzx+fb/CGKUMiZ9FYrcPw9/T6PnPotKcffdN3IhiDXQ/t1lvBC6Zb5
FkV6Im3RvdM/+lmLuckd8CxSgHL3TBSNouatpu2yMXdK+1NvRdr6maLNPoBrapfC3u5iqAXnZIeV
NGIL3az0LpmOzOJdWGnGOiw6JLw/fLN3IiiGeDFBURQRz68kTsFYXaEqBFA2SXtSTY7vorzVbFrI
lb6maiPM/gMO9qt5YFxQD8uWaBP29NEFoT7DKrr9J/MCn2ZIHPaEzWBjdxAadX0IEypRkU6tXN4k
UmDOlnzuiiSGN+3KjtBbI+zPzFIe2Ea1YdjcfSqtMOtIPIsdlZ4Stv5yu/sElE/gGbtdefUSyjIt
LL/O6qjMtyh5vxPeVwO8BZWBVvYehKiCFOeyWeWLbkLULD7e2kaxuYbpee/rRao3uZ/oXtYLJalh
YowQIQTrOkRmsZgRrk2Bdgz/G2tO/PAc0FTQqGfCmFJVyS6l9kS+dDRfi0MTZuKvi7AzFQQhZ3ZI
QjB9Ls4G48N3x4pfDrhJiClwto9MI6S8c9sseIpyLmYnVmQUczwyE/v4jgNfC5TqtkRrYaPeG9Tx
ZSleBP4ZHXTAYMF0tN9nYA4SO8YJ0Lpp/TGMmUxvLINFNhPGr+yAescj9YhQLDsjGwYuXX1sy9Tl
iq8H+4HZiW+D6725zBu64pyX4WtnuwEmpAC26LsDIW/N7RELUbVKBtuJWOBj34/tPE+ymW0rjvH0
L8rZhf3mrM4m1rAVgaWG6He2Thsjfo8XHaoeuAVTZU9/zEW6+rIuKQj11DAmQSHO4WBqLaabgpAP
m6exz4aR7zr2xt+G4T0QqKgmEX6GkP2tIgOUTXI/ZgKyR9zJ7RL3fM3vS8Esxa+BVPQ1oj9gpYp5
TURRwNeA5VC/P2WzgRxRzjFhyCIyi1653tje3a+294RMmk/6mXud6FywN5b9t2qVYgW2pYwWMSIw
k6N7a23aq2ZakOo08U+tBDOeEacrqWsjxLS3ws3M0eP8coIGvJhox2Ws6zxmmNZaPkcmc9un+Ssr
U9tUvDGzza6frWtVpJ6oOgLYzriomW0p6C0+Ew/2YL3G2gXmbqIfTv9fVKboYiKhETOYeb/4qQ5W
X7/i5A0zmTFZTNubofuZ3mbXApfca/BmWTua5h7kqf31RJpOx1KKewC3nOdMNgTurW+NyzuUL+FF
7H6mzP330b7gbLPYA7MqRLaqhtMQA4zkuBAsYlKmnS1TSjGH6PWv1zsYE6gz+tnsmc0hdsGJyYNL
G/FZFTJl67W7gMP5TfHJPOuQTBvNCVo1O6/b3DqJJBZLb4G6AT/P0aDQXuZPX2x1ueGWTvwuBSBD
qhuVFtWT04+b/R01ViU4bhmkOiUIAtrDaVe6DU6v5xrPvDJopXJSsuV5MB1z6CT8J4p2h91X32Yq
JdW1azHzu4/hrN40OuNbbEDlFrgGBm6PYPJelGSjTypA97AURYR9ABN3PtPxvNSkETfcb9CAUArd
z+lR3nMOsubvj7soDIlukiQqI/s+zp5ay3nK9aTmcvpKB6G74pnQASMfwVu/JENCOMG/1nSGC0R0
Gu8g5cVE8mZJzivfaR+CtISI8xJIJqiIq6bRPczI537D6ZjnqDVAsAY9CRCkvUDxuNghhFAXYm7r
HVy9L4EBISIJw1SL/CFr06ur30RBgKXoJvehnDU/MLWungs3EkWJP1W3TqNFPwvJ6JN5e/E9/ShS
7EONVtMFW2fVvs5ewHUt0NFnj++IkJidP4xk61SjyvxHe4+NYey9ZlNsPUccMe5Vu0zen0YFkua6
2g4kshRt9UtLyu+KaZSEPaS2Xq6lbkfuOu5F58kVlBJPz6EGs3u+nBsg+DttBRq55K4gLAyoN90a
IjLc6z8LjmlbeHbz0Pna0rrXs8YkJpFFUPjDQb9J8McJjGMWIdkylnwpr3cdRRXB/3oCqihftN5z
KcgWci5dYF+sY3QFwtV+FFwn7hoIHstF7fCcB0A4wvh3xS4A7g0k13Og57KyJV8t8lvq1nKbEEDt
CVx837rqrHetAKLGGXzUOjoslKwjq3syXapyewC68y5mp9hIT3lYsPNwzF0O4IoO1xBZ3EdTnG8f
TtSazAW3DhcEq2Myd4tnGOukSuDsCrcj8rygHwzCY3sHIghylddQmYUJRIHBoyqH8bO7Ps6ltQ9E
VNJ3v/iyAmF/Vh94Fzwjo+sTvra2nD75k/wypYR+RY4r6jDjdMmi9dcp63BCIv2ygwzLDilxGXXT
Y6pS0kvCWILWAeXjmt3+YQifEc9+EZgkQpuK7d/k7VJtrB3HUqXcQ81bTY5JR6l8uTy+elPHlC44
3vIIm1ceY1DtOUs5wwzVpfIH9juvRVRRuDlIkIKPeTW5FihDUHC4z87/ea+TvZR2kbIsT6JJg8ti
Yx38n6gWVCQqT79/hNu5X8JeQJMSl9ZfQ23sWAiqQbU7d8qIgXsWqh8zxFBm1hBO0IVdANyWYRA1
Ij2m1ZJtBZpokcC4OhIAtTpdT9wR+ovwphPFsu2IiA08S4E2B1YTmStHo/eXsh/HRFnN9MoyX2xz
b8fBLXb/BlCP+sbyQB2Nf0fo7w6Tc6muYA/KdUWn4QpTjpIgGeefrwCO4CTn2cHtvBnU1mpiPMuh
df6c/V1FNMjvWRSmpPiSYN+3jvzmam96LPzYl51Dckp8A6wg4VHin5PXwUjttEJR3Dk291FDxLx+
P0BXAgE+uFOGfKpbVy9MhBx9bzLQkBanV4JxXoGYiDbDWaZdZZaHVC6LBZxKKkxxW2iwqthHmaOx
50FJerzc5qgdUeiDNlV/AN5J2RPcwfIs1B6VKBPj0blrjMlxtDGojqAmQTOkW4kwrs2BcuQNaxNf
s7TjX0Rdb5mHA+1XAC13y+QWgQXkO6wYr1Cvv12Fw7v7kscuhZU14TKvWT7RLEr9WJPjCUc72TNg
6yCpNSbi3r07NJ7C08+reMtcyqNa77L8VK4rMjYpnh+FU8MF8Oq9QtI83F5GvmZeD3B9oRR8KJcR
NQ3ovnvK1Osdx8Ms2UHzFZPg6qlYtakyVc1HkwOV/eucLnQ6/W/j0ApaX4ax3y0fcRPfZpNvWg3n
LALZDgU0N49DyjKid2S73Ar1/KLy1aWWyB9f6uE3c/cI24gfQtUF4dIUrzAvdjgAHxZ+YIB5JSeY
Tqs51DuiY8J0wFO2+lXTN3QJEFrlPYkGcF6UMJr7IG+zw73Nx/dviBccepmFbfDdanzHp3WOx/lY
2GkyzHaR6InXv1aeBzNhrt3nVUuQGTQDCA3F3ZUJsRBeOotD4yr1e9BqFJe4T2BkUrEoKx+juBjK
+VN1b+I2hu55/4XeLgXEAjdHwhM39RDPKmJOAuvKhx9/KjAv57i6Ch4NX7sldbG0kxN9Kcv7VvaV
evYlMIGi5+o6pIKdYLYrrbV7juzOCoo3DxhjvwSCSpZDse9siBnYJb+IktsqeqF9zpmCk8mifTYZ
Ehn+EKEDTrEpz8QNu6v2xdZvye4p8pA1Yu0S2aQ8OjG+URaP0D2dl0t2SjoPykO1Dfn1dmZtgh0O
369Ps5hqTRCLXIDsvXZvAk52Y2l7SD81Bxp8Nra2GXz7JNwtoN+uVhTWHCghFpTy99okgQT77eD8
Ej2kQiIYcG17JJm2HMJ5jQuZc7V7HOcaZIinqh2dOvMq1ydwnav7o6UwQHbdVm6dnJ+kYBzHOEoN
jT2N9kHZ4FJnuCTDXbs2rmvsMWOPCg+PiYd+eWNRMLtNMOotLlmiBP9u4aqpidLu5relnvzdRvt7
jKo/z8pxVuTmM/d78x0Mr9wf8xPmDyqsVzf0QTnYkkkpVAgP3xs5GWkO3VDrssBAyl/Lj81NkL6F
w2743+RfNjhu8WfTnfcOBwG2izzIz0VKpSlQokuhFOnDluc7YpI9W35rahggGfEz0+lMqnokJs9I
aqfZSnHtha5TYjztuopXS1CRoGYVw1PAn1GOYQXMxbIFhv2AQvFgEd1nonM3qGB5r66UI3UNKVue
RRCc63MmNbfYVNxybUVxpI47DFtTS1Ifm9kTPiaAdUVgBAYjabm22hps/AvhepeUobGA5Ni19ds5
rgfCKgTVmxvmsNPAyURo0xSWYrv3LMbw/J2AfPp7nTVrtE/QC6C7RUHXiGHp3dEujkUMw/GoudMR
10jU/0c4xMQUbqqyVf1cl8mQa/fM/KjfQ1nADjml+FPqZJ72mSUrqPStMpkpYX7NlrAn1gpNTUbT
ipa4N3G2lkirLslYWIWTM2/BHpLjJNyddFYdBhBD4J20JFPXF1umHLnKbAmIksEBmfakkV5BUDdR
19U25LOI2CTKUSXJfKfIwVe6r04VKZKGuJit8fijwCZ6nNsZM+a2inLeGD+xclkhcfHY97vI2YhY
6yRyxh/vrmorQ3aehCdC2h8UzH3zDSMBBbLcrbucPkm4F/WzW9C6S0VzfSlJKk2YOGZHgh4j4snt
dRY5aibzbq/ThNDvZF4dCEU1zh2rxlVw9w/lcDckld/qwHo3zFth3YD6morXIXlC1vFmC7WQvUsX
WivEfUu/BcftCtDovvhjOwIyMQPGWTodskMV5fe9MeSyfgyLcamD4PvITcB5ZLoSpnANtf9MDhNz
QSEwr4yyUj8f827XWguHIG6nqZgiCBw9LOlYThScOb7Saed+YtZtAsCct3YvJwn5UTUCPVl/yLUn
EQj5v39ZOgeuKpSDe7DiUYvCyilHzgp0aHL638wbdE+c1AwFBPJwcDGzz8032dR4woDA9snAfmtN
RecaeIp/oEUkR+RtD8wrPkQFJO5SkjcfMQOYVfD7In4tGG0KKDuYECcZv5jNThUOVS9dAQ6Nl00Y
XTFIAgSUD2qGEb6njgk3HTi3qLGLudaoe8/CAeafNWeJESV+JBgWKUCRY/a4tx7LRLa6QUEeqewR
079DmlrPwGbYhd7+gImpc9KRLwU+klYhBfkbcPfpMj8nCR1Vaxh/XUEV/uQojwopqo1+4FivUvJL
ueUBJicSg/34gDmSFh2gn2tDyfccN4WK3F7HSlsGv/fLbL72I32rQmCxBmjShtSR9zabAkGwEk+x
Jtwu8H9QE9QON5y4fjNTYR/3+0rfFa2PedmLAxPmPE7wU8M8xhQiuyeWakM6DkxpFp7E0olRp54R
IGQ6i1Z8wryL/XnHTO+CNbW5M9yvktfrUfQO71BCC20KriIk92ReRTwapIRCxhL1lxASvdKdP8hq
saIf1tnZf1sXgaj7JNfZpPW5ExvZpAnQwAwd09avJlZ/0DhzV0kNUcsYIZY8gYVm8f2kNRAjc+5K
guMLc0QxbDPwyAuw/zID+sMZKtWdVYpA5GFfdAZmiDaVvZtfA2Sl9pFg2vmC80D51dO2f3ave8x6
7Gy5Biuf7JKbRn4iHBI4mOiidBCngP9Q3KC7of8BjN7g+ujlN8Kj3dgY9NVhaA4kHSgFdwk4Q1CM
qum7nNtd2mgrj/jwTG13N/mEs7qCdIx+boGTg0adgFV/DttZe0b+LbAIGu8DUzz1NNvTyWYKcejz
d5z2lSTQ8x0cBcBnyA84Q5bkpYutfFdMR4zuLemWeKxiapT73TIMqpSyIrw6ILVteV6f06kxB2ow
pJYsu1h2sCUfQsAhYGDoMVCsPCL8WDtw95busMBsu8Yf3/qWHION46jHz5kdjlyNNDRDd/kXIleV
1LmAlfsKL2EaUxqe9dK7lioIJ0vn3NEcHg/35tIvgFnNuDAK6a24sZ6Uzw4Uko05+T4Fcp0qPhw4
ZfhD2dAtSfqBHxyiqoMp2aTHKJ7/aZ0Kt6cCqvWQ0OqZ0zpFm7W6K+eR7cUARazlAKwPakwsDXjP
HwY7vvmbU2UT6Mj9eFrJ9ewEmViYHdXtyXxXs5aR+06TyemsaF4bl3iAwyY70/tU6pDimotKm7jp
s/nC8Bmj8+pvqo1NaR8dAdc+s0RcUTixQcvW7ArL7GntN+H1B/Y1q32nfeCLIyo0FBweBZPGhS+I
iLr1W67FHJ7TrSXL1qp1uO1qMIDxpIscrMa9kR7B3DIz0IL9dvr98la7tM0JafW9OARKaw5Li+Ca
kEQSwc+DKozLIDcbO5EqvNsHcCugB99q5Kis3/MPH6XvZT+o02/KClpd0zbsQUaWvB6r4ScoNZVc
whx/959wWCaXXSYe08zZ+moyh4Gu48mi0HVtvqhBesF67K2ko8SVnl+IrmKTL53/3PlpDp0ahgSO
84mSPLAmVxkNvODzOzGdZmvED0nWQgN/PYnKcNOZnMrmfJRuX143qZiLmp5rDNiUSS8ZClZQNhfm
F3TL04cw1IlOYZBMrhs9GTkkN9p2FJ9ZD3cYkook2yzkYhLLNLpd6XRka3bkDwe0kFHrwHFg01pl
3Yh5r9wIRuhzihlcoAecAQeYGfg+CE8spqPMl74gwqlGs1uXRWoDP1aKDIBr/PNKHyyHUwfDiapy
k4W+qp3bE8DRbhaKkZbL/AnyVy0NgsBTCAtmaA9ZJbN5753ifvKYQbx1IONY3DB1DHh+EIMqAPwh
971PcIRgDv0PFb6ouXy47GdUMCDVGUUhdJDQDeijl77ED5ff2C1CeM9B+PFALCAL+FEQDqQm2dja
25mEOGlOtdn3iThxo3WGn16Sge/3ff2dy0C8gVPiX40cn4yUd6vQuAc/pbB05ZaPA/UbWtgbeWmr
vCO+Xx3TpoXwbe65EW6iVO39ezshU5d9iY4RGYhwDa6hKJs2VPuwP2edQTffthNuOKAcTAk+JuQ/
k01E3leuVy3Lk6x8BIdxW9C+Uu9GHiS0VJ/VWtvY1IVwXffTn9srpuR86wsN5bTV4hnJwKwF4zEV
nyVLoOf3NUaTv2kbku9+TNV4US8tIir7LmzsQY+/ZvNsti80bGSXisC//b3hAc04CdEvINCY85Y7
gjJ58htFq1Rl3WELimKJMZXK2dRrPjx+byOugyeT38v7Veip6DVZtIN/F0kjgwVW5X0l/J+XEcEL
rqTbkMnpHTjlbyEviXUOEfAYVsOB+8tm0GlR5cof7Rvv54amdb8Nlt7Kq3ZNGON/Z4l63N3E7Nhz
Fspf2wJ5y7qhyVUnTUCx7oEt86QN1OrSlyJE5aj/cB9YjYvjKEVzTwFjqhIEucfs1Ud0dwX9o+Rx
GWZA8fqP3PFReXxRxb5oJnEaDhfGy68cDzpIMuzpkjJTEVtFD/UE+8ACMYN6eQJ1dRy72ECfvZT4
R5OONtdS9z0gHozh8dZ8WdnYHvm3DixqwfmFvqc/djo3TFzno8cc887+I5Af5+0kW7QRMvriUrkE
8I/g4wqgdIyOpAgxsE6Hztr4ljQQYlDrme9I+wolb+LknxO8ByC6jM0ijWTLSF0lR5C4IS2EwhMG
XBdarCTYXKnxg1UV52CtUtZz+JuHRPvpinvEbzzBGDDdcfaWt4RQ0eW1P4aMnjJ6hxQH7P2qcY1B
QIfZO2UZ16R3r5qW0F7lR8KVfvxb9uMqo8R65ndbii86ETBpeHkxIdD1CObwTRMOnq3VaVh7Imxu
PN+3IYmdCgFSX5x7jDG2whjW+veAo9TLrQdfxhjQUDID4C8UYGS2LBgvffwBnr8ZzGwj+n56Qydw
tMA3yQU3DM6QS/Hr56qI34yzY0nf+FHGnKtjbw6wslgfTzQwpTL+jrnpjQ4Cdk7NogjWr/2y6nJc
BFZ5gq1olMekaJ2CfQDwHW0yYrVXe3wboPYYMjwTZ/NGlwAcyipqzpk0O3G8es2116we9XwfdJkR
x/JigWsvXGdVQHxk0Mt9HsDebpDrOBe0s0R7dXjoT0DkoHu/h73nyFG9Jk7/wX4OLi1jfHCoKci4
5ok8Htf8SoiFxna3RxD1XocY2XrUuyBXcxyQ/6Gl7Bd4W+CaY/nwBLg6eO4T6kthks533yxCkv4Q
GZDDh8QGjo4SN4vP19KrxNfLXmSniZuIIkNT0xK6MKZ9UctmXemGSz+VugaWrZQtJVZHeA0FPrUV
w7IC2EDLODzW8QflR3GeT7pekEkdRCAiTK3rNGVwxM7bLM8OiatgMnVCv43YPWI76l5RqyoRcikk
zMhZAegWmtcvFdO+itJaLr4kmu+g3gAzIvKD5jVEWn0Ugmm3YMic5bqesdZS6K0RWaupgYVrRay9
0s2x2AAhySQBNdCrizMR6OYAX/8XAFnF/8Km+VzmIWNt8bGrumqxacmdvyWH0PSBcKd83QomYfcM
OvC6TFbQN6yX7DEyMaac7AvNetdGUUIDQOU/DnYyWdakbPeOQ2Bp7yw2e5zDP7K2EvIoMthOCd0a
GgN1yphFAsoWIbPwQNn0/qMGPv8bOI/CJdyPY25mg1oCgyxneuWCT/jXu6cARBB94gT2TlI83uZm
06LO2w0zdD2adXGDGI7uM+QorhUL2mCX3gYhFZ8b519XVa8RQ3REL/fnMuykJisnYFR76wnzAlU9
bc+TuOq8gJGE7Jl7CgpY8dtIWiki7Mo5RdetDG31qktttNGZGr+88iHg2SZwP5ryYE3xuwjFzXU1
TIZZl03yVOfI7ei1MpqzVbG5tlTXszxOuycv5RgkTgpMByFwX9yAjcBV+PBHAiKCUHO6YaKNx8QX
2sL5mh72h3mqA0kedBFl5Z6dhzV5gN48KsPGS8G4vYIeXI4n8eCbzSQ8mb4YW/lbgqFKtkE7vseF
VV/vxfgUt48hU0zDken7bausb2iY0T2jleLsUgkVRpY1IYEUo7jakQWZEFEGpV6ToG5Z6HN2hTso
yTp5eGkraYqKW7qk7R9Vs0gr8D+QE2KFviwJYgGMVrrvM8njy5PLIFgros/Ku5oW3KAIdbgC/Fny
bDgSLDwqZqh0h4A7pkyU6VxArAv6YHZEZp6EmtV7Oa0PPdQ4K90Ltz2+Vmc47LqDW5PnOf3r/LwK
IPXgsJXY5ymj6pGOQt1eyvdZEBasPXdTsGp7zmAc9sB9gu5yJbzE8vazFcAtp+ctZCccnQK08h6/
EnaD5O2pdKF0upFMkIjnHCz+YrfdASHy6yB+BkrrIYRD10MTZ8L8wCQ8T2Unz/jfTbxtHqCOyG4r
NYuGTdEAzFIXrxfy4h6cGhgoxreYkYNbU++0megEt3Wr4nr0BPr3NtA0gb2NM6kqkhtrRLalYFGH
cDQ8z7nUbslIsxskSBMfmmqD1IEYw96vWEm1nhLQdj10ib9Afh7+hLCNL0UqG0iIR9FuzVSDD2c3
RR5mJCTOUXvpBhwEptcWHQG9JuMx5cRavSkiPYmHwgiEj4MDsY0fTPQSobMWzwYWTDNiC+m0aiZf
cf2XhJS78PTkOZmp21zA2ZuKvN2ZVlPuk4ThZL0xfd1O5Qsv0QNHJqflwVnYQTpinJpIZQOkZdpN
z80pjqdH3jMl775YRiIpN/J8/ksnGeATysN9Rg1+VbyMf4QMO5Gu8yBBNlDIuuDiZqZl93vAdn+V
mHuw8Sg43tTsyljntD230kqBD0ZtRnpfXfOB4ZxyF7Fm8+70p5SbdnGSQpj2sS3Xpnu8uL2LI723
wXxE2eC5X6NdNB72Z6mG7D4VASqWGw+dpQXc9t/jlYvYVY9UploBOaRVD6fQVzrbJz45vtzibTkx
KfoUfFkxlD4qet3QwPF00H40LrfobzURMDbnFbAj+Ga+uq/D6aq1p4Irus2bRsfxEnxaKFiSoX5e
eP7fqsLPm4AUy2/om3fk6LCdGUkJWhV04JHKIyO/S+4AQQUtduBEDZFOeELmKCwDFEDsykIb7KyK
vAfZwiyezOHraQjEWsKNB0G2cahQELkDtgkPnZHG27cz8KlAAyk0QdfDBdiXoTap0EITKcwAtE3q
kfgNAEfeVn5t22tJ0wAcyiTzOdX3iKXMqQ630Jqgtl3TQWq4mA+V9gr+p8nzbYtx/wrChhajwY5Z
bNeL3A6K41aoJA1TLkDuZxanT5ADs+XXqYp9hGLb+6HkUlujnFVUharjuz6brWNFqAYzGarxG22o
OLvsko897bq7MGrGnktekQA/eJIxhrm89YNB5bFFFWzbip1L4uZcuUNA5P1qaQs6h5jz7crxq0yH
Dvx9Ma5Ia7hEQBUGO9BIbrcv6NFoT4pdxhlKa/raJl0F/3+DODyAya9tJX+T/0dK4/3YyG8AjF8A
nYHWutyk4pt143EANx99tjLjfgtltZif09kpMKlBR+8/KdEgbc8CiFVXS6pz6U1581BwH8qxJRk4
4orcWvKnIIh/cdc9TE4HF2p7HTGwic+jzJomEJ5FX3LHOR6yAZBwqh0FDlOGhv06XJ85q9ASf6BZ
I98MHEtZfEFREO445SGcFgq+rl+AYMcVUO+LePW39oEAPrzOl8Xn6YAnZ6ST/2UUcreU9Sy8TAcP
IjxRGlzvEaBCKS1VxAb0x1lm75XIdcgTNj2dhk3j2ogU2HpGjgXm6wLceWiBv7+v5iV+ngDpNzbC
8Nw4nKye60CxtuzfelY5UrSFJDbVz7q9YuXvdRhH3KBsKq5/31Kxfe5H15ThSD1KU8fYI8q+eIIs
k39okCmy361FLT5KIIMAKeaNaA96c8HWc4abNlg6F7eZadi/MOK3GXA2msieay+An7pIy/+RN7Sc
ik7xa9GxlJ09sSxauErHA9ochDA2c6SA9anQHAp4/bwe9dEXIV5PoRcnWFYjJh2PbT6kU8aiOO9r
VXwTY6b2DNjNTxKn9hvGSXc6hb5UniLSEpU09RLZB5RHt1K/F+H8k+tVLaxY8CWne1iV4gGbnvUr
Y0uPr52j384QBRHwUMTyzgdXQAqmi+wDrG9uch/TQsu04vKYr/xpcGqNxJMxS089gymVZgNmJ+TE
fDtoeKECaIiA81enQewgbOB1V0klyT5cU+zqslxjrWhXAvJkWgyoMahqMudIVrTJlIryB2FSVoBV
gDOF31PndeKEDDkN+K6IWTo1bD8w82kH2w6eJeHZV0zmNYbPyJu+DgGnieqTsEJVsUp135udGODn
WM2j/wItWYyAOcNV1mFKk6/la3uHS8A379HzGhk0YZYpjSjWJXM27va7u1+Et79TA07vMniL+pvH
K9zgrF8wixbbLPJbKMK3smONLfx1DEs8fnJ7qkkwGFHabRFwiIRJlhpR76zWoMC9LwgMtMvxZ7EB
ttYAEOYIy+wy7kcjIMXREcB3bkCXsYpdukzy6QhNOkFIbaGxiRWPBgkg+UWgs4hrGsLhPFXoBsq+
DN6HVfYbA7YjYNk0FM5cznIc+4hGFBHG9Hk7AgfQWPFawX8uP41fwpUaFOxW+pWttcIHNyfo9jmi
t4LGr0p28mi5a+iYH8nzLMXhcbE5MTZiTT4gQC+uIpMe7Cpi983k6Uoqi1rVCz6t9VJNQV7uNof6
X4J6PD+HNxGsaKWBQaQ2BpST/eb3enIHidrfjl292de08IwdEbKPTaberBiwfhZDtmuO8S8zGy5K
4HUoeVyFPOYvfHwnixYnj9MFWwuxJcWMuxLq0JWsEbm1DF+mIgoyUSBYXlnP81an13TtOLeIcG3q
cRrQuWm/0N1EG8OjzU5xQxswGyf3Swf8yvD1fk/AONXxS7MzXs7hHQEKg7cM+2uUgt5USxySCxNg
aGJGHdKdpcRUpCxsbNq2ZxfGZpY4C4eYKhDlYU0oZmpe/FkKuGfzvQ7dOOCZMeHkHWqx2iwj3Fis
iEZXQYi1Ok0jrQNjUEx1/7euDkkzWYMRKqchz4kw+EdNcqMWOdsxexQwxB2f8B1tzL8Aiu9mYfCu
gA7YtW8Bspus1brWNRAJqF5nTaRkQwyk+RI4Q4dMA+BdXKtsY1ws9RLzYCheTPJtJ0g5ghjKIfHL
vDY5R5Dusili2wrtNEeA6Tf2nzRVIUC4OWg8HY3vZCk/03j+AEPRf4bV+5d71F2eDpa+32UQuc0T
9UQocqRc2w/OpK3TpIA3Ps9mOhZHIomGBTxa6EwahGd6YXZ3uoIlPVrjn31sPErrYJNrcIWkT6ZV
Iud/H48YlVEMJIm1oAiDQVxkZTLyqbWzjc/dwhdVVRqoUhg5BCI8Hi2Ita6MXZJ+yLiGSjQSh3wF
MSb2x4PLiSxXU5vmdcguRR02XvgD9IxRd8VLOQ59YiQ+4p8cZE1fp+ZZljjNL7AbxRVV4IXfj4/T
AccerOPqUQjkb6SKNC0v5BP3+h4nWf/vNZa7h45kik5HAPIBYoh9JGEDDYtjgbFB1wRiVN7fDA6f
WZIqDI0dJbgw2RyyHFGipCaeiTGnhj4KyVbamf2QlnfNl9hoGk2Yv1LuDsl8tDHVJsfQiaozCSkd
c1ELIOVHNMb3Afibja40/4fPnJa3hU6ab1dVLdvsQ13k6TKEpq/+re10PT2+khzACLRudew/9zWb
ZzHmunJJhgPXoEEfrDhNgXngBUCtGZ2LUq2rrD9p8M0+iuwcTwjkjwld6TCaIpJHdzplkVmSbv74
zrbsvsWnlKTg5+8FZRq7M/XSGhXnpY2sdkK6PbH7eWdhJUj7jTgysBiW0sdjzXW1UMpyEJz81iwS
CIWk/dy3nCDf0wGcVY2N4odPhn/tYU2CuS5Gm8EpA6c5JJqtia6g+72KmEegoIMPqSug8l1jwNO2
zG3uQo2LejLiOnkwpf7SnKta+h8ecn0gEX10Gg8ZHLlUMIPWAEPiFcPykEUj4j4EGjxxOfqb11zt
0TGDux8+aFhNkYPrtPksRBaBW6YooRpACCJhO0BnsdYeyutOZlY3NG3AyaJc6cvPqxWst39i+zvM
bKlyv+U86JhF5RiaL+r55wuQy+5ZjH3yB/WrspuVkFWCfw0T+zC/QfLQ/kCFeHXbx4Wx5sAtYFeB
IKaK3HUQqsSDTpm5tOq9R7sP9Tn45MRSFD8AfocDJMuC0CNvag/FkAh01X20VYTyr9dmW4cFlPXc
P9Hlk3M6LHbyl5rF50t9AqIDFFhF6jGtM16tJC/bW/RUW/7ZeYEtLgPtkYv9Wn9ttsw2N+EVxgPk
dUoj0zMTtZ3Sr3lREMuyiXT8ww0haw8v7X3vyaYlSbwbcaXWfjHnGAQlOZuWoy6t6+yCRdjDM8f0
HG97w1BuDjVBDKdINlhWMU8PjiMYr8Yqmsnpx1odgk2M//9yPNDZj7OEBVLMUi2o0yu1XJobSTY5
OJJQtEqPMxJlwRsIA0qLhUZ8gRP581nivRs8G6QpgGqLy0fnyJCVlgDJfjQyRVRxIJmXaTriW8Jz
MjopB1c8YaPO+FvDVscXRqS9yst9li0ZecI/UZeldJYBGrs9ScxW2ZWFO1o0kMcjmNW6SWSKSy51
bFfK+LUCy3pJbChYoQ6VvouV3JlzprEFEJs7L5rw+uukU+fZao9mEJsyqrIOjH8YP8SOnmR8/o5b
rCLgX7cYmWHZaVt78Xo4UX9e/+7+C+yehZrEz6Ki9v/tN7/FRYPKaP/unQV//qcZ3WGsUIhrfB1j
Z85fdWfssQvA2N9/TsAGov1ZGqRQQXvklmzQUWhReCtFcIB90HMshleyQaY6wln8tpNWrB4bFy+n
4FokwE4fNDxpxtEoQyi/FcIKyxPY+EM1m2dwnyvNYfQ0Tyu5sEopQjdNFnTpKkxrxoUgGfLbHGbu
B7A88/nBrt568CGPsJpWsU/qCtMZrKsjMkcKgkGPcUmCp6YNpo/HGqoBxSeo+K6VCS81YHpb2UwT
waW3df0C8ODUBfdaVjylJ1LiqqNI/EnPEEsrg2IRNPj7yFI+l4tOWxe4VIRK0/428hP3l19FsdAB
TwshZ9ozEFTNRpvGLO1z/oFUvVJwZOH+hRGo4jpIO0cIDfvTPFbTGoa9Ix+ERnslL9siYer6o3zM
e3cB1366+n7tr5VrR8uBohGnAG5gT2ZR5kiraXc8pczG+2VkercVT6BgJHa6ypn4rbuWIA0Dx5Lj
7ogWhIoGtAOes96AuN3VXlPjo1S449EH9O1w5AxidRRgy+d3j1wkswJEOS1TID9z+nzIjF2KxbFR
+Jr68Nr8W7C6ar/ctKseee8hgYzwsdNqal9/mKFZgiqbNID+KjdVvsw6Ip6nhKYiCgAbLEuzqoz2
rIgBhb0Cmn+Nf4uz9nss8IBFMBcmY4/blL3h02RHBo51tw3jekMqSQ2O4F0x9fZfljqX0VAIlwVn
1+icEfYqLgTHGVXbSFfjzqRoz/hYgTaxUBBDiUwCnBOZB/nFwhQvvbpaQc8ZRhkairUMGpmXBeIF
RbULPC9olLT6A24G+sytkz5pKTJal/W9qtkKPX7mR3s/dBlUTuK4xfs395v0bucAdF9ojBRIUxPu
fR/cBxUscNTil0cDiWZoeKva8bBpIKMvZjs6Mbo0L2APwQ+LLJ9dCi+Ic58EABRHDMPmeVUBy4Xc
sIurghd3PpWtDPUpfHSIrRxZjx4zZZTAAYPMz5yFQHz3VOElnBJYorGbROUrwIAGImuAIC21owB4
u9pXapVyOYnxzboYoHeYB279HqnWO64TlJJUpKyxeUcjKm0xfd8kS+cpC5NK98PXK0QXWvKDjpK5
ey/1669vyXTNiZhYBjgbiObb3hsffRnrNenCk8RSlXbeUvQUEk0rlWbKQa6Zs3lFpmhWL5/K7xFa
w6Phsey9tT3LmkQT82nwBvJnjjpUYQvsbi1lP8SCfr0u4xLaY6XLXu1IcovgA6rvhqKMVi834m7C
Q2efBP7iWuOQfsqdgjQUt9nClVA5TyS3T4CHbFDDtW8Q7yAKA+qfxp8GFltwreLYahsb1avE1ylr
UFO7Orfc0haWXtQ0MIioh1AjxO/orwVabyXeFvU7YQdz0+gTNIbaidWMJGGMi6wG24IvkuA/TpWL
rOIiKrePnvG4vzK6dgb+e803gsNifGIhbyNUBAh8ag4MsTubtc+5XhLKk3uT3z3vTpSVUJPAtbAe
Vj9ZCdIv1P6o272XfA9Q2k6rY+9VYu04E8oOvTg6c3YQ72COH1GWf7O9eeBsmF2EMHfnvnPfGtM/
J9PCPuLhLZrIvuAIQdddc8lGthyRFS2GVcUHDIUAsPUv6adzKEni24g59VurM6R3jRuWUuOaj8hl
vvGqKkAhvUwlCfZH8hp6N31v1+uxpTVMljT4s/uyR3lD1SuslH/7hXK6EOwiZT/9KTOHNufQWtsW
lUS/QTnXIQWAha08dCVSLV0H+GYik3DVT9pr37hTP7FZG6cFknKSnbBcLfRMtsBQvNxAzLjJIhCW
BIgk+cPwznl4Ig9VJ7D6UHGfZfLU9b+RSOCPUm9fCQRtQBHhrvyK1DpyaSUw6NiBCbyvaUDAevVy
kW4V8xpgM6ZYnOntE2P/t4YPSKNY2ZWtcJLZL//czvWW052lBUQRIR6CLHn5inNY6TtMQEkXaByA
zRRQOPI1u400HZ25qKh8YOcuyXE9y8DkvEgz/7NdtMZMAbIOjW2SO78O9sMsMPmkMCp4IDHoqVCe
NMGYTUe/vzOPNQZTxzoQZzhrQYEMDjYgvyT3VlXQxF5pLLDXupXIYH+Ezja8liUXpzw5o6kEG8FK
g0XAudWSfG8hb1BV6JfW40n2VQICEzpuN5SyyEF4I1GHPMIdYoMPL7pn3JYh8fAj651tf1kuo3t8
tWxqK1/u6I858wwQZI1RUEf7b4yklZbOmgiEtQ+JtdD7jhb47Q7ktVVTCrwFI18gKV8OcJWB3QxL
EkWfjOKOmjya0h/R/eiXf1s1+sTmkfIChRroV00KNPdBLUQzy/2NZEl3JcGiiMCS4Lmg7Zhrt5dO
7YEjvukZUffHE3Dbo6hJCs9HOrUHGuEgv5Y0lzIW3yDzuhWvsbuusAIbMb+dQDepg3ZscX4UTzNM
XXCG/DZDdcvsgdadTjhNDQcvyGNgT58T21dLwEAL5He1l2aRetxrrmeMD1Z3Q/Im0Furk9ZxljDg
yoxbN0HcYaSriT7TkliVlj/NYekqLhOboqZ9OCWbqdo6G+aUtsTE/TyCnFuVJy1CgvuMPDhyX34m
MAjwxIibtxHhB1/NaizHCoKEqPcnSFtnl00xpmrE4/YsatavqdSP87TPytHOExPMYxHCjtEuKncA
s0IS2CIj/JDO/WU3vR4LjSke9jvdZTZmA4/8IgJOpJZvybOQo0yazVpHa/bMA37Ex/Qq8ZpyUk+e
q1bZNvgGXbDH9JR/QHnCwjBwD+S4uLrbI17uCGHxtIwLvGQJsBSu9j0vuyioh3kcbr9KG+fkpukz
We8JSOf1uVJDTlVWfQHblpBtc4TT4B8AwARz+Q+D1KLaT+NAfvVjIvD/NmpYU8Kq93cY66GBshX9
XAUJCM8JwWExXA4P33tv0LHmT89tTQQEcyG6hP75srI7c6/2J5JUkfZQB1sN+pXvmUsprO4WtOkp
HXTcqq3oZqgXbj4TCUqiJ1+4ZeIxb76Sb09p9roIWqm9bBWqj8N7LIo6gC12jzGk3a6k7XRyPG0B
hU0Jv1YtnOa4Zh+g4/4eEBqR2X9lRgdAG0/Y5sE1Cfpa3hFvvzCzEfbyhOhCvuyPsWrg65IET+98
bhfK1NuFpJa6FcRm2yMjQcRm003gma8p+EU0qk5X2xCEMR1LH0uXNXZ9MbpEURruxET3gijgHXL3
DQViwpEv/hbyBJvxArg0Mi1VVEAqG4SVeRm74UfBVGsHMkGlSKvMxTgKQGc9pezxa5M2LBmdsvYT
1Uu3o2hOKqOraMD/pfUiytaR5uXCv5O2YaFmBy+v+q5f61vRL902M/Ivb+kxWuyTWSY9L+WY7bR8
eEOnZAqaTzeWmVTQ4KG8u0yTIKhEPoCN6JnS9K7zW4ntYLr6WnZeACrYNWlwHPlaybRNBIWAdm1x
kRn5Ic5V4AO8nRd0Ne1ssx0HI4qVUrfDhqhi7PiQ84nU1uivdjMFNyHkFZU0wkKSmm1gTCEr8Myl
jdtahkbiLfsKsrUVlE37hBubGjrGTl04zrdUIS9q72vQXBn1U9P3wcJ4U320vdP1Em7DdlGyaChW
CmXjeb0z62FazrnfMYyc00lDv9SSkxOfqP6mRHYzvC57PxCWN3YXD07XHdp6VrswtoNc2fAlw6JI
TDDqQhXG87RShjbQP7XnsmIS2iD9IY3mNJa/ecL7fxBkMTRS9P16xo53nNRpj9sThfE/Q5cPQL4H
iWAVyXbszU6haghF/C2yiQPOcpTbS9SqsdWPCdF9/qkmXcFh+H0Ra9ku523rCgzAzH8aXYbaTwLG
9WSdlWtSP3lEiAPShWNUlfae00SUk4H1nkrbA4kliMwTL2NGrhLB1Fo1jniolN579MnEAfdOyJNy
jBJ54MK6K1VFm52rPrcCZmRm9HngTRmKqtHf9oS4PsyzcDurfatLuSmnvt6YhgcMlTZjXFKJizVu
TSoXrrZ3qbVOKFCdmoRQniaVcBbimvrwx8lZTwX2rD5ETAATHJSQpvq1mevLdOz8khKre/v2uzqn
52lmYlPw07THdTx5XwSxaZhH6Ft1pQHEc0OqutwfEWBvD+lABMo/tWhcH2i681OoPipGPWJnjSMN
8CCG5+YmMr0v0b99TmDAyI41sjLsfHVX/dwTkfciKRBYf9Y+eJNhfDFN0SwbwOFgHZj23Kfygbg4
a2+CNshzUENUc/n6QlyZXPdUd1hPNejQPlyqgdhE3FaP3CPLSRrn+JtYCbWT1gnmomxOS5Erpnd8
TT149Q+kA6SLQkSPvOs04aIAmJkas63FNd9zfP2Pihp6PC3ZDmHy5rYh9e/DMlWzkZnii7a1csj0
cwzT6gAy7wSTK7w4UIAohdgcehB9nonmU/1WWHwXguxlHU0qVI1Rw8FRGcHALwpDLssrncjnYlL+
Kjv8bbodSqxy32isas2pWhmPTUFAXHqieMjfYMMs/m/B97xP1ApJTcLt4YYXYLOnIXy0sTAEgUBz
gj75rxF/eGpgZo5dJA/naJrjl1qjMSpxsylUwfd/2qMOO8pMaaF7HUAl3wpvLn/9PHoh/D3eWvtl
L8NdApAVmSWm9EQhNPaEVWUFqh9HVZJADDMBFcsyd1tmmy1b003pCbOu/jHXhHqfDOePsz6OS3nu
cbCpU2t0iI/F2RPajIk0weqfBrBzBO/rdC+jtzU6XOrcuFkjGuW8SIXvP8uM/cbohZxjoKL7c6jA
Gff3S2M2RYYbbM+iGjUebkI56hb9rlPnTmJ5CLUzO9LcW3Imu+PrAtQd7LHdqmOsTHmdfpi3/OXT
WP37XUYi2G7lM6t11Fp/ekWycvc8CeGTC6tvyFcst+Jc/dT72EemiIHN+R872di4ummbTuCj/PPR
1u7LkXif6iLvL3q1rQjMdANiLpByQs7yClLEZI+iLZ3SGo9epJbG9tBYT/SRDwP8wTGM8mL4JRRy
F8/B3ATC0JGjAiDisbhiwe15QMd6gFKnhk/5slBW6fFUIQhRubpHkR+WL2UD2ZBTKlGhguPN4tiB
I6yU/4+VpK/zITX8Rwj0gqpDdv8pEzcwL2woZSTn3Er/n9eSJBtxKwhrBI6Qz3wZIbxKErTg5KWy
FAHxDcKKImwu02LWhr8Y9+relp/EcEQkb4TlHdYZpC2/5TpiFVK7OjqXwY3CQvNBfHYpKZ+GskR7
mY3p6S/5CCrX5LfAx42A8DNffw9cMlG0e4HodrifsXH97j6Ts5/zqF73ZBLJeWOi7y+zY0RWeacO
KFUirpnB4MWvWvu3nhACd0LLTH6Bd99VLA2K+Paof3igmvIjCtahJBcPXTnRBcrid6nRqsX0HnS7
XT3kpXGqa4Uw9jPmiC777ksp3evNSVqQaowv7ELzIz5Gm7wBcjHma5E+Ud9DlLh9TpA7/t07C/Lz
X/ewATt1fz/cKbKsCCaKQVi7GoCx2hKX3IzspR/G0u6BcTMdwM3kaXfT4lq2AmBc+VP++xVdMKnX
L2IRubinz7x7T5joBOcBJfskEKOBwYtUnD1SeBkILHCqcdMeIWOhNnrVNUsO/YWl/RjYxRXnvozE
O+4fEikv5LtRuw1RuJVup3phqMiShUtBUus30oA6UrhSyj0mXrwcwjof1aCrzaNjo9VL1dYA1ziv
GpQVQ/jgzVIwulu1VvbkYWa9KULdPAbrArPfuPAlfGkvw29VP299vIv8xNLYpEYAeosSLmkinkI4
980ZwFA1XGmtvrxaxp+gmhQeLPEReaZUvQZfF7FfSER/36psUcWqcPccJwhAufB1g2Q2XtZ63BkJ
dmlqyHm/gRWqi8EKlLjxbnB5QtzaUsTTmKN1wX6Ox2YoysY+NFPrYpjsmER6GpGUF422M6cCEZjO
JZOrtovwRon9dB8WXdBpjf++2VqweXTxHYvMhdZNI6sqGv1kI7MFHWHGYSLuCcrk+ZZonNsV1Sue
KU24Qq4pEHtwDaLSSU2o/uVwpf2YALWDPCBf0/PUyLHzKnetcJ36bbZSXtukZcIXw+G+Us6FkkDa
8xfvgBGpHrLUIYm9XpusD7rmfh9Cv9G5CkX3qifhaOKMQK4WBQQoz0LvDnDDDXWQcRPzdysFTYbZ
QYOjht0clfg1C7pkbajTuW7WxuqC/ls+y5Vu87GUIcYuQjckyNpWnrJV1TvrJ0aSt5cqgtjSYfDi
xGfIn95th2YoIQrZ/7PDdW0LkJ9OoIIj6XrTQA56kSCaImeONy/5U3XdEToCLp365MaGKrLovn60
SGdXD1/Hjggcy3zZmWA1Yy5QQMznFxj0dDY/TIZZBTCCFvHC6pbZdIBuDLBON6tbsZHT7Z+uiXdG
au1GraL+K0LB1rjF+SrAc1hiG8o+M057WtLWak8PTddZCh33i0XuKutZADX9JzWBR1llNxMezBOy
7EHL8jH/IJkIGalUH53a5y0e2P2MLoUjj6NnwNRJave0BO84HL0MDANHQjerl9p51nh+lD6i0dTm
D4xosWnyQL+AIe/R2zgs+BFhRJOiZ8Jg8GEORwV0bwMzIMFx4EpiCcJrKVC/a5sqxesXe49o3mN6
Jha5g6p699JBwvqCPWGDgooQXstAcg+EX1POOHUyUYW34TvmGx4WmbyMpQgYYkkRRnwhlaAHrkrq
FWvGObkmlCKtTDx3QAbrg0eLO21fSBGuISm0JF8r5WsdzhFTXBL7bdylgUnjK0ahOA7aSayuDF62
k/v12l0wHKkSNilDFbCYkyF4EMpx34Bs5aFO8qfuuOM+JJ/CK7XWR0CHQvKB+3CBJHzwu10PXj16
np3zKsKMzaiaPKUSPs4tNY7USkcz3Vak8+KvuLOAPbL8OIEZmNjTF1k6ByJkatqAB0dySMf6DCUl
HqY7YHJ88CqVOW3CBgQZbIhPPME0gcogNG814WDbNxJkPc1uIm3Eebp/o1Xzb6BDqGUieQN6ce0v
sZ1kXH3AElO5hPNPeL6AM0Xho7/KiXtqI91d5BQaMY/zI1kzc+cOTjeLG7eu8mlL/eOevIATAJw4
V0P6+/Yq4Ij5dkMDUAGkCW9iPUcYiII4KY0jIDq+BOtPT8mF/4duyfRonPAJqWaY+dwURTeZs6br
Q6E6dfbmYl3BzvlRTYVByOVQLFOWNm+rOLopTtIV5YJeMCps86dQE/8PqwlBUqWidXMFO/JfWl/W
Xb2Squqf1hWdsXSHJrHlLuIWQ3ZOXs/355k2E3KtEnLB4JwmIGGeeVQAVdEdTzflgu6ei37UqwwZ
cXM+ffwrjXKZ2ZyaDCJT2EAKVxdhB2+Big7CEk3g5v0ajIqZMeNbI2Uxm0d9KAsddqomO9Nkidgj
x0YZQOSl1hFxpB+sNGbHDMCShjfxsTEwhWrGRuCHxLxzx1CqYoXrD6G4jD8IueWAFStqoi2qC8Vi
dgpwRme2K4XNMFfhwKs+7t3LYPpJG9NOO079tfLUyUgqCh7JQXSyUq6Zw+Th7cRdm7p348wFyEfD
7G4XqVjXELgq3c/d7eaIRg4ojEhn+M6+6M5HRG4BSRfv1m1BiDAx2NeGAZe5KNguQRm0QFkNGaAr
dzibRQLTMBcTrGnxdqSNgxd530GgXYbSgESyNBUumKPkln2/6sqsZcQ8KJSt3BYZQbarHQeuU05x
YzE/Rsoy5hvbdnJvMpigkxYZw0FFbqkbNnhTtx3sHs35Y4FPjAGT7wNgFWxFrw2ygYPrBaCOeuHt
/cRSPf6rj/f1npPlYTboCAV5Nawu6GRrWH6bWRexiHGoNMnalDfAkFU6w93KjsaUtuOHkwEHwpOi
RvgTIw62kTktPDu26QziTMm2avod8xb3tlO6hjQaMngW1XzkAmmrd5f9RU1LXEPx6sjgedfWwZuz
uxfh6sl7RFmOXYfkaAlEOXb9viMIs2rRjskZfem4LXa4Nt/ngPSZcn2HKGNoxhBjuSDkFLvvwB5Y
WXzPGXz4sTfS4mQAk4YVk3iho8iuHRK7bUoPJCl7SQPz1voO0CKgOyTYt3n9qmrv15YHkkfBeqYc
QkhMro2toysHWYYpNbl09ihfX7UVQEVAS9yxperfFzBXbHMLFvf3CfoWlrPgC6qn/bWD/n6jQ8FB
3AL+ymgPeUa6ARjto4VYC64aU8L5A0UXg5vTfVBdtgAATzEtCNdtNWG0FrYh/Q74bdcBOJ35eWJA
Bja7wFIa3NXK+d877LTAY0UG7Ic16b74vlZ7nErPs1gqO94KqMqz05lHTIdd+b0hYklw+ut0+Qcn
YDTe1g1ZGW7saMZaxlzBmQX0MiqRtfP8c+faPA/VdC1eYMZyakkBlrZldgoJTXoQzsdOHa833aU3
8kbUjPPIiUQJb90cE94I4iuxmBoD2OkfKwyBiWfWvTDBWIuyeLu4WhriMYd0nfBDC/nQZzd1FkOf
mkx0sNaYKDqBTlYj3dGOKvVVniuDbWvFCOmaweHX4p6WEk3aprcaMa61uthqftoxxsy955XY4R/Z
Z/ZBtlIoiWJBJAkD+jtXZq10pwTFkEE2ssW77VI0sYqOukGE2NGB9Qx8KJ6Gh09UWXEecU7O7MLu
6uEGCoh9n0HYvXeTnTw1bIsCQz5yVKNocxPDG2rQw2jyfN0+R3BRavE+wRPzz0vzcfYPGDQgV2E+
zRo/Gbx2lw6VaOW6FTJa8fIP4XjtlVGR5hkyY8xLaMc9luf+5nfdPVf5qPsS+ZXmfRV0TVP3qtIC
noP/aRF7O+s0bD++Vx0UZ9dmIf277F7hFaYHxt7z6oYOJeWsoUthF7xgmTpZ4u1b29RORFc32zXv
5yBKZoj7Qf0a7iVZkZgZcQpJEGaCdzHraYKQU+S9/KNQLG+pb84rESfMLOdJMpwSK8WAHhe3pOU5
YS0QaGQP5ST7U71TvHm5dl8EC2a5N/JJdOdtx9tMeP6z4Qpo1fR3AMZZr7ITG68DQGH6lOGl47E9
hPk9Z4P7brfvM7oSO4ockgRYUXXK3u0DMjrhtPKJShkgv0H0fOlQIOSU1f2BToV2nzNUwE9Pymc3
AH6F7qUNswDxxv3VLS7vvCjBcQaZJyIV+pcwigrPFRoBOpC4Zjlg/exDra+RQTbLaJdKEtJ6nAfq
rg+CciamI3pOJZqO/fHP/abgdqYN5B8cZevRFvlqGm9jBPwHt2t6J1jQ+O6s4kYpbaYWnXId88o/
5X378XRi/ucKAZNiAsf981IbmFgl0qO5AxFvf+AWJQ1PMWtXHBvljN5au0d3COXekx2sYcgieM2U
0uFo+GDXfnAA0x+AsIDPzvO/3lk/a3PqFcB05cwJ1XF8Za4hlBwaMuY/4g+KZiuhVMfvk6EZu/bQ
GnnIaErWPk+Y5WL96aVMMe5+br3J9alpM7vIJqaSus+aTY8nX9rHPAQKI6924/RVG60c6k7NWicT
3riebQXhFpubDOzLf1eHNRmF5k+962GPhFa7lbCzGGAYuwA/lSQd1uKzZH+SQ57U4iediGxYdr4v
+kNnbXNYdsiG/Ftuc3r9qK1K59JzzcVpQu11i7Rx6GeMSc0nt/PcT7HooOb56rXOd6fGyF3itqvS
KELrBtInLzfVmev7IycvGUGECfc4V1i2Lu3yZIIOfPGBOD3hC7yUcF3bZYGXlOy8dzuFCOZ9A/Sv
Q/nNJxp4WsO9xnRoImTCVA0o/CLT0ylCML5FM4ZR8CVtSyF4nFC4RwGhYO8uiKHGfWK24fWufqU9
VU584XAeVvQeD/VmwOmwa0L/Q7Aw1+uVbvuwspemX/adSXqFPA5RGpYlHKXIyWSdSQeG9QO5ToZ8
GKB9j1vfb6GpIYOJlpkrEB3zFsRuAjLcF5udMDuOU+rtKmy7vGv+yrQSQBQzrQAvEDHaXqrRh92P
iZiDS5gnl4RfEiEyhDOlC8siBivUS4bvThpOu6Pg1MH+avrmVSidzwUYNJPBRr02bSNKKVf01iUL
NmIf+LvuGLw5ncKSoWDgoLFxTng7K9Jvuvrulhz9Z51PjbpNnNZqRitKjvNgXaQoBSgaks7HQ/73
5Bbd2lHwPOwfkJWp3zGHW/y6Q6OiPJXMp3IPV5RayzF6bISxtllOhiX8cv4vfvyUoJ3LRUFOe2j0
Z7dbB5oqUXBtdDVBkYfcIu0Gw+RbTnbdeEDv3UsHdvrZtvTeRIWSRLt/rEaDQc/xvbE97neU2gv5
PB3y2znsee2uPd288LetQqBbwoYa4W3OQvHk9y+VqGYQ1OVXzaWZjCDP+c8FlaAkAIa9cmU88Cyn
kEM0ZLLBG09SyemSd6qhqgdt4EgWbrgLcBRql6P+CF0eC6cbcsBaDVC3SLViCjtb9rnGue3L6o6J
RwXB2rO32i/Y35eBrcDFEsjcHaZyKW5q8uokTHkB180bk8jllupZtfq1SAiEZAtmXxWDpHDNXNA3
737weuNBqcmEdrqkpdrvUJKeRH8M7pJ5NcqEoWTqm6BTL7INGPqeFCe2L527o1v/MTkWaHpFwdTJ
Y1FW8bKXRgCpN2HMNpPsr2K3eV0Pr9ZjEal3Vtgy7WvrW6h/mgz+IwKEIpBDM2I5rLEIJ99iCbKO
i7NuRV2uyoymuf4AuFPn3I7gAGSjUFFBIsiqE/l6RCHKbg0wpu2ayE4tvMZhFJhTwvYQGVOFQNj2
x5FmmaRIA6+zQYvOAYpuFr51GqHGXUD/vr60XkQArDqn746m0u5/XKW/7G7wq50fs7N1X9sL06MI
O482O58EUdRODGTvAFstPJJyqmWpyxVMgqJFuxf8j8bzWQFWKX12O2x7A9mjqkv9oqyRRg/Gban8
FOGaRZbgtjE1NeRtMGJECnUtQgIB9lgkY0NkBY06zeoz8H7l5hqSYvS1i0UhdHzcV+r4XROdpNwA
k//mwWMm7MWIWXdwF2ys43/EoHkeVXf2ktsKDD2opdJjsM3ziykluMO+O2wwXFJSkyTD1eILSeDu
7w8TCEh73/UjP3EHV3i7u5OVQOTHjMq8jwYjEMDdfn5Q0b2lVraD5hNnkKTMP1dMwK4uCwfTSVUf
uQ/c10kfMkYoHoqhO5tmb2/XGUyB/N4krBdmz0lL7HVqBFpD4+jN8yCPGaAEf2mff8BNTJPJi+AD
x7gWKNucZkZ2A1C4K+ckMCrQ+6qoTQlGXmeGlXZXHzKOhI83ZKNlg1BW4qEDSOiXO1g4CBqZsmLU
mMQ+AOA0K3rTkLMurR79Mcc/yA0sdHD4UE9RxpAIEvHihNfUceG/3gnGS9TmO5ZSvk7lVf5Clr4O
fQYW+4rBdn8PtmA2Xq6D5abahS5uQCpJ/GpTifdnkzsxM//n8+18Pzt10vq32BCdbYw921Vs9H/J
AQKYd3uEu1WBI1LVem0+j7f67G31rq+I6syDhd+wRtuwp79m+27yr4DrqHDURUfwwip8g3s9MrtY
BRoFNK6GOjwvPzgC8k6e+munyKubJaTEML89Nw/4siH+lmgFCNPVXsNRboYh9fb/wx7R/BLxibii
/xNArQax7jrEveKwnS83Y3PP62CvxH8KNWp/weuro8miHbTRpdqmjwq8EP9IF+wnDPDxauCBXIoQ
1c1yeRlJjYEf1/J5L8QJu0wkgyQY1IzaKVT2UiNULBfFNjHEbSG/sIZLwrf+jq5QYGydAcDq1TDC
eAagxFvuNXhNlxVlhic3abhxRalBuO0m/MI/cMi+w6uzzgse8w9+nYGxyJW2ZCEBfNU5ugBXYXrf
k//Nk1woblwNu66PfLWHuL72s4ws1WWkot9zs4Lu4ROYLw13EckrcLdAEgLWCf7bBUbBpswygt5/
2y7dPGUUJqW/zTeB/KSoJB6FLCHGsjYcSnkOnv+gnrV63crqHN2QWgdAOSBnpdkmDvm2xofMGuCV
lmI0AD7cr7u8pe/kza5XcCRPcrk8svZru3WogNL46Iy6cbkCFGEizxxqmhxH3aToyd1kwzyqM9/9
q+YoiqnjS88KRfIcFeXub9DHmE1cLWtrOxXTrgIOnkrQJmf+pNPOL5oWi0cZ799++GsHC8eYSYEt
kRXL6X3CTQAmGf6Ugl/xQTcC0tbYTjMGJ8i56F8jMGIuRoGxwHz5bVuEZ5eouE1G9DzyzIHCe9uI
WJ8HUyqCi+jhyiXGTsebmesGo9+T0pVmV8tMfIjnzYRUN5/TPgk5Ec+2kL9hWYxGdOWvHwxfczgl
IcRFnwsKzNzpVoF5Fb0mfV5Zf0G5GaxEWv5yZTsoQnD73NeCOQUYhIXlna6RsneyQg2IofdugUEb
j7AzFrr3aKhKpumErnDUSokNliHZPRuYyeoiSFe6jaNCmJEXe5WDWeJeKhK6zVJlj7+Sub+/lY3F
n9ejjoKDPh3QztKNI0AK1j34vRGtevKhZyY8GiHEmz2x4czSqli5TU74uX1anXOQmNYXZ6Cb5aGP
Q7cJ8wUIpmOEjq4D3Nbf372L9aLgs3HvvPQcpSQ133QZ615maMFNnSrC/wDpLGFX/bmIm+c2OzZg
GfuzTLdS7h7AZIDvz+LpntPw80myoMtKk698c1L1gSCJPghhyt18tNqnyl4mvTHoGIW243z4rVf6
VveDDhfs9hcJ8TmyzH4JH0VjKYtSmIZmy0Si6NE5JoaheZ3+QVZrwuIMgfJ+oMzuNy5UDHq1q0zj
dHPzoG2nGrO+taAzxlbyho2cvX62wuUK1niSzAXqxG4Q6OtsNC9COtoBco2ac0BR5YfGFq7nJMca
t7oLtf3gCZ2IUaPeFFllH7gii6RNybUTukwXbmMnQRbxv1ZbXvpPJR6PiqxwnBkH+LDu4icoB/M8
s8Ty4RTxcQAMtOTeynTHm/6fVsCFF2Giy1MY0Jr66XAOSjoiPnKzUjM08Iu7IbUEwqADhvk2J/Ah
ca5wfUH7lNyZebd7WVJOSqrnw5IGj7Yks4yBFyd0IUGbZkRoAwoRP5SPUPHnq1aVcfkFEbGZStgs
aXYd9SdirJNCa6Udbpd+Gz2eq/NrRAGGZTyw1EBek7X89LuI2sTE+b7lMbAGej2k4kD4lxmt28ME
mHT60UZEwP0u1LolE8ogDezDUvihzEpXOESq7Af6W53VykyeglppWK4eMJmDPJhPU0OP86iYTYNm
jh6IBdrVYrSO2l1NExYul305T9KQK6JsDtJOOWu4og2QyML7h13STOUSG5fmW0GwyYnTPHkHBjT5
FsMv9Bblgd6Ms9BW3gZFbBFcfutiS+N2wAqk1kPczy3rUSkWf1AYZBZUwu7TsAg4d3vsc8z0wH2d
pWNok7hAwGGtDz/NPGENY2YKz9kddzahfEoJdxi+sRUx/8EdEdcKWtH8v2jO73EY7XsvRJXCOgUf
kMn4K9Mr+yk9aa7AJTJgbFJ7Lk1au2riMKpoa57a3/NiiO3WhZbjZ9bM0zJlnKj6dJuy1sWL1UFS
l7Gvr6tvMx2SMNPpUrJf/8x1tnFV4FFIly8zJcfakV7VGYpzXhX1RWkDLPuyP44HTDa+sCL83Wsf
KHDew5ynAs5QXpnSaQ/mE98VtWlT+Gg6IX9ikSiLV6pFARkmt3cGJAbeQwRCUktxQvcuEAiaDAda
LUigZA+R4lDjoEDM6rYMCX+iW050c3xDLPfz0azKE5YwiD7PAhF46tk1jPfcij28tdL/v4JzZejU
G5P6g6i5S+OjBIzjIV3ibHgT55FF4sl0W8A9g+okXb7Ye7PpgAyz/l2kRvqWJf89UXNId/kDrM1p
xNXVS11Oq0+OPnp4DaR5077kBnnVD8UlFQin1qHSK+N53CX98R9mFQlHFN+Q17m6NrUty+q7y/VS
mXCzN4wPPUSQIlqHzXGS33mqizbv7MEJ1WKB8njRckzZXYguDUZzyvz7DFhuy/cjxDmdbBPq/bUZ
j3vOGzV2X3XBN/W1z49pikp8cc0IoGTMR17zDIu5i/qAI0W9RHMAxogcSgsWNW8xV8HXGnX5IoOR
hdoueyhP2rUngquzwE6LH71BmL47gPHWARt9TRMmDhMaSmPJPFwwbi4xEt6gX3K2XsyZXNy3e0fR
lbETScUliAfc8126tyfew4MWspwfQhlUPBxn9nqD8q7AiHXFunVviLT+TyWHW+5nCbsfzW/GtAX1
SqaxxfuO+zJyBi6/tJMWGa3/7h5VRNtm0zgDe1rSBLxawzdc0fMhZHbMZ8LvQJu8JhOt94hseFIr
Xn2Uke1pnwiviBvKytOjiyulTI0GUiXurOScS1r3Sdajb7bQQsHd/wJNy26XZuCD/19NFAFcu8Ab
h7qHLNprBtF7wdV6ug8aSNrKe2LAHty6eV7g7MUNHcFnbKainGDIFudqG3hnx42xhiQw8cCVGnK3
TJQZQSbb202KKOeJs3x1SBXAbBdP1LBDxgEz7CbI07L976LqBYxkTE0tBvCJSTsEuhpZbEvxZcM/
x38j7CG5QGYvg4C+OhTlHcMbDOf2kiyfBhWknenNtTJ2uItW57pMArvJFkdplIt8S5XOAcRVhOr4
pPMM/Ss9whci+GftOWV6iwfQKC3XhLuhFmGMfbhXNZMdvuM4sUr3Y/F0Gex/8UxG42gnCxaMvCV7
4JpIMx2RsTYCXxMBN4LZ3jWo8c95wyRC2lQ6fGNPy4FX8hlyuhE5lbAZGox8UiPZu2hch+XLiQsW
NOZ8om3LvzSZ2IYdf/Zvg+0ic9ZWqt3luJvnh8Zh/LX5FcmiAg0chALvG0K9EHT1uDvxUQJ7Ja/o
2u+yCBteaVref1gwEj2LGCCMI1bqufmXut8dH2Nc8VleaMvIl4PqNsIjPNvk9YEYa+CdTj/ERyG1
1XuZiDg+Q4YdJvyI7tNZTw8lsGBnm1U2kEhlJKGEdrtlLiB14lgiuEqtK/JYSpxoQc6RJONzNtb3
xMbUl0kFAl68nUs1b1/T79tCAEIEdk6popNArL4ENPnyjo6Fj7/uGL7yAr5f1+RVIDELWNpAUATf
uDeThK7R1/6MFIGmgK+lEt+ddw7vXB0lY3BT5/jtLKiRC2qAJKguCciQdyR/F+HhujtY+IJwkhtv
lUOwSHC5FnLxgh0uqri3IgRsVn2cRp0IENQTe0LCsokg+j000kKsOU7nvqRLsEz6QOAH/Dq/eUxE
1IQ4/zz2B8U9fNApIj9oWJMJoOH+AWhZoMSeDBmJYNPEvSURtp3uu75YzRtWeWTITPbbLY2/Ijc4
oxO6YPKaWXeLwzTWwngHxkth4NhPcCLEo3YSa/YiUlfpGhxHpR6kOKT/GuX6yEBFsnGtChqBuoSx
N8VNWwEeFywlzXyLzcUYAmUMZ03DbbSFpPUMLS+jX+dn66lnT/ohIjfZX6VJoqeiDtGKkeNOWPb6
qC3MAW43mtYIWQM71wKOEjBF4FB4c809hixYJF+E8fKzl+G+wIr39hc0NhOdS7TIZbMpj2iuZo/1
zo/wjt9rAOXCMLLdSNHdS6IT1EgbrUm4CZcHuJdYG5gi9QHuAWQNYDKRjW8FxDKM52aAkXjPJcKm
a+W5T3jmWgYOUxkUbgZABBRmuDm0VCxdtsn1kvKov7XqJteZAgowGCC53ghAiLe70w3BCF3ppA/w
rNj/qgOJlzuqCUw0TES61UZnthbyYR98GKe5R/1x6gq5pmSeQP8PbV1UTdUqllmqDz+K45DNsr1v
FhDeDX44RNHylFhTAblpgJB6CcB6pFjIhlKihAkhK798B+7c8QDg7qgUHEJaxBguIuL8fhbpi9WA
LC2O+CPtCq8bX94PBuyZK/KMqFLa5QVXdWCSyE49Cn/ivXEHM/8mOxyoy0AZXYnAqFA8haQNSNFn
kYKTAdD/eE3tZt1ZOCGyPPvdHv0sjSroXsoYufVybfUQW9NpcG9BiJ029Idr87yLIXihvb5RMuQ9
+wfBeAjdthbCecoVd7G+3zzmdPp6452ZxEtR3qti06mlsYchk4oqzt5do6+espQZToPVHj2Jgnn1
AnnCFdEaOAUl+Izwh6f4yL8Sd/TtP1wv94wXnt2HYqdnHJZUHfv6ANl3QjA/WmON5aVevR7gelHm
rXSHNstrdFl7+R7HV8hbza02kzhYJet8qhy/SfR0/gwILd8Qj4hxLbBO0CgrX4Bmlbo5c6rRAWix
xN7HqpP7BmMzVtqpsOf4z+LpcgNqKXY01G090DgNSQZJ3l0wKopFlsOzFzdalFPypHTIneulaVUj
1x03lIYpaPVyMiraf2ns3xtjTgG7elXDV5EKo04jKcold4IbNY4/yApAHjuXYxXWZzMm8eCvTem2
rROIoubPqGb5s1tRiK3rE7rA2iZd6i2PoOYzzczrTmFaMPfSKc/6buY+LjSXS0BtO1IsLPQT/pkN
Pjg+nSBkDWLCAxPuht2rL5FhzYSqDe65w+26tfZSYSk4J7AdhgT0X74UQaxYLM5HgplhHnp0G2g/
5E+1ECcCLJwPy+NfjHYFp5z91fdSxlN+AC4NLMGy5aNcTtJT+kBzcMfYj68JNsAkv0ikfiDejE7P
dZG05srdJ/lUbmg3sjs5ac2Tu8QkiIhYwKY0G9z6XIyAKSEd/AM94223Pmvm3iWNybCcMma1jDf5
w571WeOXYmWhWmt+QXibY+pSeFmrWL00V+aPgn2lEBlBgfQwbdjUL+ySdV5nkHr6VbBe8QLPYmeJ
ylyGdxvXMsz3RZzUuRNGoIst18wAt2un73BbTS4y3izejOKaKhV5GDzyk84d4LUKQVnn475BOrC9
wu9oMAWs89ktN74e0gttZQpzGy3LAALLv3ARujVGMuXeIufSsZuBbWn6u7p9H5Ir2F8P1YZ7wN1M
aDDhYx4ZjKOwLUaRyvG0GRwuhowGMbfJihFqzm4L9Fnlv7bK8/N3vc5cqbx34XSN+w+uQdD21brp
7UqFd3uJPWpBefytfaI3naIZzKPOYjYf4+UywdE7Wx3MDBwcEmVt1e6xldRo2SdBTxF6OH/VDye4
H7zL2bLk0Ei81khqpEb65BN+yNRhjC5uu5FmLdSB7KsNgp/cEMQP5Sr04EVDPhzC62HW9XNkKZqH
IbIecIL0vtTqLD8E562C72CYj8QOW2dzWnqvh6h8hEGi//V/ZGU33M/sd9RuGj3nl3mwfNg7mF5B
qLffZebcrgDHv/URIsbDK3PnMLtDp0+o+BRVDhv4r9SqvJiGV4vJSiwTsGtfeOaIq+0Wuvlrfip9
vvI4m5ve5gaGCPHZHMUdCkcxF4CPZ6OdwfPZ1G/f18VN6jIbM9PNhhSeHica52HJoaPCpcGE7APF
rExnbqK/n/uVtyniSLmxv3J+2yW8uLxjrrhcwJDSg2nINjV5symGPxx3r9PpDxmaEvyF7e5YZNEP
pTnzdD8PpjtFngCoPPENG1A851J6HWnle0ZE79g1ircFYA/gSoWGvawti3Hp/gzzK2ZwxeZDH4xi
ftkbVWLj+9nG6SQepV8im1rMj+0Izb/zfZ0xhBdZKfD63ZD4CF5MOJCP9T3R6qFyWgULqvEqbXDY
lMQdwkPkuKQnhvMfaNgQ482cG0buTQR5U83rCLRX93Ob4Ca442nF1sUUr4Lh+PV5dx7tzEZqgd7d
sXeBJKBc2jtxaHk+UiAHo4Jw7TNBo4sEv1bHQ1bAUhBsqx8WKXw9KTq9jT7aKQvWcPTcZFT8nMkD
owKUHSbljfDDnyUyk5qSnLDLeaBdpiDUda0PBXzYOpbTTgBCcGYuKR/DpQRjUEiVEMlNsFcCwKup
tBBZCHKqk+OJspy2l8d4/LJmPXU7pMF4AnZyEe62mO2RFtfHH9uRvcsfP7BSv/j20i+HUxDgkeP2
jAmMQGq9KFs20BIeIKPZSObjNwx3UN+Sfp4LMM4r4lEXt+74ZEfEdny58V5yifTs2RjU2qsZRu3U
rG6k9MOtmPvVdbye4tcyeSddl9B8DKsVOZJLuNprcIm7tEvXozC/XTgcdmoEcR0gf4ZVoFvBhigG
PQYrE7wtsEDc6xfY4pfzNadtsS/XohRg5/MVcyD5XjM3WqXkwBF3s5FayDBiyAG+dsU7sOH/2qvt
IWYiffdKUBmqtSI5J278AZZGx23oQ5oY69avIrvvsIu6uElQOVJPPCledTyCQ8Wo/GBwT/wPuTQZ
u+9ZBz8vIL0FnYaJpzm/768QdWiMinhGX0TqYOFmJ3EKZepGAOOHbZqzhmcrTX6zX5VlRYOADA1T
gR50Gvcr9883rNE1x/fZL1PJG3UvOGKFIGX69CtEKppyxqyXKhudbeeKe+0scX74qS0yBbFKzzeY
Q/wnKNnBpz09XJmAfcwBzqxZUoJxO6x8yxuLR3RcFHh3BDaxctTORV4AXbU6t2CJpyLTmZE+qtkP
QI/oyMzajpV7DgrbyO6nanSFb4g70EpdRTVqSbokoN/eCCIu6hgbk277v596cO6aSZClNzzevqig
6+2vhywJGRHJUGUFjUfD5wwhVpfzwjRGCYqCZmh0soq8gPTBj+r2inybnAKOup0S0A/uP6ZHM+Hj
csvwmTYme8fj2XWq4UphuSBGKb7DjO1t6oyJjk4ibwSl7Kve/c72jdIedcldO04ktGSND73lmS/P
WLXtcqbxNJIomV9axqO5Pr6XETsT7wibvda9it873o6JVTupq4PmuP0Sbju6JQeXUNP0UIcqc1A4
A3Pt4zxTPlJN2oVR8fmAQmtIZvIyn0NDV6MWkoNpTkCS0feE4ol6t2LgMda5b3+2Ev6dJnR2pApJ
irWvBGrFCWpeQlj4J6ZTZWjEFcFQTx4Uzh2DYllzjpQ9BcUYcHrtyP7vjejJrOJdf6iOzOB3wBX3
CyNuYXkfZimNTu12t7Upd2Y14+2u0CbOOCWMKqccU0Wt2RXEsTJGOaREoCWasQTcUaLmCzY0oQCW
f/RZ4jrKMhzxGmV2BzrdZpckalGWjZJ4/GptvK8k50C+DslMrp73VXcXJavbtNs0g+YvdqZ2cW2I
EWTZO6ObhNKC5hQhU/Q7kDUarWwFeA5CicNTKuef1dXExOuyJJgDnuv01vOTFcRFolcokKlsz5K7
r2bVRb7wid1k+MihB4gfpzQhr7NwjPRsQRwUwQzP7oUU0wLxuB1cG+aTIQ8NqC0AUC/701ietgQS
6RPrxWcWLpyCrFltCtuX7lXdBfB6UG3rT11DnTSeKTADqSVme/VZ8C/fZFcOo3iW37aMdaqrvGXJ
5GhzdRh1DWH62b+v5r3/RqYLOK4vOG7qhbLyBUeZQu8lzaGkVGGuA68p/cxVhn/PyXFeOIz9p3rI
0hFAhbebRj85Z9Ejc1PWYQAHFR4ygbh3GmQyzg/f2WbXswl33uP5ofpYeK2cUXHeWvTQxw2DL7IB
NZfUEKplqDc0RUmxMfBXlNkHYBWRhSTSn2eXm4UNpbW8ITrjPL2QDZ+mgF+M77/00N89JgvmrIXY
0mzIhtBJ505SNjMWaMt2g/lAQzjH5e0/6YZgNYoZqpBkJWIPTOWnseZZ8Szll3pKlNu3Ymd/Ot8B
P+9FJTD5X1fFwag7g979HcGDMIlZgtCvjlDXmJU9OV1YVpbUMMp2g041BS+UQa+pQkoFajXTpqs0
67dwG9fMSZyTnev5wm2hHry6z4Ahbq4X2VO7Pui0VIiXKdcOcrvo1xdcD0ObhWyhNy8B1bE6GlBI
W7QAO5iSvXMnfz5u6h1Kpp5ZJcMpmrea9bI/N6fIeokWCwukw1BFXnyyIRvaJOHLAOmrKlmW078B
RebAl2N5tU7m3Vjk9E3vrRZzBcVf+/dQs7uY8l+WgCDBLKeLx1hY0w5toTi5fvWVkTGuRiWgwneV
MHwm8/7hhxqgXaQO1O1swjJ8dXP0AaYrz9GURNJ8dRlP9yDgYWIcetqV1EJ6icVYQQcRJkSucDOY
Ickj+I82iwFkMZdURPKZl/Yrk5mkIVXQ818LbdvmjXKPtdqmEwtigxEqFcCZ5H9Tp5VJPO+pUDSV
QYQW01U4oZKc23RPPQgfcPYi3f1LD/4HvTzjHqMZztMV8PjaL2pROoGdnjYnjZo55bhEfcoKE3zN
kVGgAkFyJlSTqHNCZeAz3KZFG2RuMYWpGCm7bN+NCCL8Q1hJ2N4qcyBtqIcwrtQln/YT+EWrOLBY
r4Ko4mBKFLYhkXs3Dn4cWARrJqmYVfw0HjLrPcWkq0kdNKYSEoPZ+LbyQB1cR+JJ5rOC9NI0uOdn
HjsPlw4MmVL8ukJUNMvOhETN5vq25bempfrhSvCH+/aBLRQTHvQk5hfYtPvQgmO2O9Tx4M0Hgyg4
9qxPBRYi/qfQVOyAvrOOxr1PE/gD79aE9G6peH6S9VVD2QRDqG//ty5t+73FeUbkGzf/SIeqawxI
HHNj+8LjEf1RH9Vm4ndI7D8mElVjxrmG6yfPiilLXRUMf11nfxsxRNej7T30o2KfVjYbgiW01fl6
oVf7FGzcPIiC/UIySsEsgVH2RdFGk2t9Dj9eDvIdTM8YFyaAJRRM0/RrbeiY+llGV++VvtL4s51I
Va6aMSZsbiDEfz0SVU4U+FZnq+dx/Loa1d77slSW39r7HGHrOJZ3GflDnwdIBfzj5lAP3cpHuN2b
AiI/1IgJrDVlWplWcSQL+GoEbGmKw3VkTrU/yufRZhSQO8OWYwgztd0nrPfMnc0ra8a5HrhVKf2e
/1mfEIn7V1YdrVsbQZo9tn/urL0JJlew2VG/aI6YQmxbti8Rp/zMqXU8k/OgNaIizyjtWeAEBLC+
kMrmENgMYZk5GXjcP2BOpsQk8Bdj7XFIp1LBBLhOEh+08Te1O8/63X+Fxe6oX0wYAN17ChHrrd0b
Ifhnbsw801+knFEacawwGaJcCCYkg5JBHYdkiLzaxf2o33Dl3bkHpGGmaqZpqdxC9vD4aDmIFsQV
dJPZpqd6H6lLsQHeGoTHDjugWavQ479MrqVIedZMi/5bPoxEg8ZqOSw+DHIduxZqZORXTtsmMllu
J1eZaGqSLePaGuxenz+tx+WnZzy10AVkynCf3Nn9EmKOoB77VzVj4GaWUyF4LDqbk0BOyEvoPkfb
0oeU35VNLDOX5B15OMmkSU45MVlFW9SRzxYQPlYdivF8JwA+OBPAYbcG6uX1GKRdjNWfbOULfXM9
tLg/RU5v/sIr1sPZtUhKP9EHzaEbG+ELWcxuD8KxZcMkdWt+j1uc+bEfOgOyOx/tkEl8bB1PqbiG
haiGpS9eMst+WTymEzS1/Zuc6TiI5RiGAQpwK7/DuacecUe8fxmskmNxNEZoXBCu0igTPZS0PCE3
h5yCu3NNI6+fxQsiExUzef+H4zvqovw9vmBaptDFUcsayj2ubzkoKtCHUMJHkPg8+YvPguSkSL9y
zyGcQGRwXFsJVoqd/3mmttnItyCjgKgIBeL+DOOGrVlqcImOTkg/yEeVQCnjDKPyFxIPzH+gPT5u
921GdXuR6Yjm3IczbT8e+O//FBcFUmtwdaomcsKz/4dZCcj2gHsuH/M6kGtrI0NrO07pE3TDzEii
mmjyElp5NavZngHxHqol6CxIwn0oCtKvbX7HErhY1c1WNY02ylnvMQp3pdU3mrjJH0C+rcx70W3I
Kmwi6ziavuG8j2zPNSmzqPfkygZsjgo0c83w1UgDsjlhcBkgiRy38y4VKEWaKTzxgLvjiWFjFUBX
7pTp1cOM0CclGvb4Am+kTBjLXHrCvBQ5/7heHEsc/+oqAB20P8+nGleUTWuX9LrlWW86dYvCrYKu
J4ov6mbBHaVF3VcuG+eF6gRoJTQSl3objlZWWZuffpFrcbpi6oY+JNrPAGK32YPnWRdM1Efo2J/a
dTDDdpGqaQynpajKmPKYI6QIRs45HNzi3YxQvCfNpKSjflnBNstLwfN05+68U3yZaNmuztx+fHYN
PqXrp0MKxfMr0KwnCpGKANQoTEEfSVKPUZNMfPeSEzDxTnUMFKlNEz8+pnwVIdTEp4jjBE1jNi04
DigBooXcD9DPa0Bz5JMG/TPfb9KX1KHI8Tjfw/4pKq0WVl/kj/cy7iQ8C0RzMYruY+Gm1Fp3QkWu
dnAoKSAAD3bmBc1xEPjf/UaGIVvuytOPaRBciHiMY9AgTHlZtCTHrF+/S/nctwbjxTx3yEumxQ5c
oGjmxlz5JN/5oNKNiW2ptPQKIIUZR3wgxBNPp4s/rDbcom84B6qXIDTx/htsxufx8sS5ukdmyOSs
Yfm/jwhoPyjsTPAcnmMEN8dYs2T0CXae+dJ/1GPKZpOvbg+WV1WpegDozxIC2JtJi1IBr4rTXwN/
btynMZL3G4uUATzdLwXFlUpVmgOJhKuQ0JNW39cjXSeXwI6J60CQU+iY59Pwu67zNHRSQBxQWwhL
M+oxVqnRTHjagTGxFSo0O2M+flpmbrSBB1NxMO8MhwJJWlvCSskTdSTJ7cutvWccV4xTsFwcXngH
1Z1GxYvIaVE3Lfs+eClnnjybuW5Oc3G9QM09Z/qMpmNHOw3JoF+WVlKAfiSV+JhViRAeG4b6C1BJ
H6Q8KAVv35dS6x0o2VjG463xtvbFS1JWgHpnJX81IXeH1kuLIRF/4kkfPRiywUf6+gMz76V53YlC
7pXIQ0Vs7QylpIPonkWeap0NNmu2j1i+vXnrKldt/m8CBwUuyh0iH+wXmivVBFbGB9JllSQMJHHE
h/7T05kzxP47Gs6Kzg7YrKTe+5u0ncGqIUJWK7CaBuR6cpIuNEaheebNuoF3/Y6U0BthHOhk9lwC
trFL+Khg0KclOwFngMPNDPHBPxaFhQ2CayBZVigWAxTjTKoPK6IXmqVsADssEWBpW1sty08NZTR2
RnK9RFlZvmHbzsmVvks1oolBgQQuIYSwG6KPPBiMIPfoLDhLeh9OfT0pzGJi2oW2Jsvno7RpF17t
ounpbeeHEJIYhd9QROi0WxIJl41Q4PIljlfPb906ysJY1VEEHMVKZhCNUTXOJfpCgq+rKEPF5NQf
qg52KdtYE9e5rnKJephsbAwzLm2ktOAUZAx5U8Vx9+z7hbM2wf4Q+V0bNvSw0f1StNzOqC4ikuC+
WrWG+MVrXSZ1IgqgOEpMV5Z6MgYaozJXdlKsYcEo6g+ngeNkWSuEV+bbtgZr4xnnXoGht22sgwCr
e2UIOSe3aHrI0P4CEk4Hj7hPa6iA8wTqBEp+vCghWHkoncQvgI264AULXvgMAhNfErjQhbDJgeFa
H7cjnFFAlI1q6yMXwR9+0zOWyx9moSi4t/W+nXOdI3kuHjjm6NMmHcA4F21so+Mk/d7UnclYt10j
tRXUDWPsWluBwo8YrjOa8npZNmLDxFTyI62Avy/g9u+Z/7DF/2rDb3hugdp+3EcFWOtDWAU6Qi/m
U8EV3GLMWflhg5/W+PCBIjk4hSFnxBIAicSgsfPpMjhq8Bic5D6SnfEsO4Kfn38j34TZVBcxwrm9
+vSgAmTynQVa0wRk1KUul8Z2Uxm8LUbARN5dcq9k0SR/pg8LBqHcD2r/ggdV5a9h3F1BdNkxjCXR
rAGkCah9k0iw6Vhg9pLSnZbikCzJqG4CbvE/dlWNiAj+03hWgZQmhqswpO/afIu2b6LTNTkfNekW
JaDLKccIawDsS6ajVzB+KZtTDXj3B6aTNSpDPtW0xL+/7qM9fkVHVvlIHBciM+wQ53eXhF2DlD8B
EJcy6sVcopS0lpNLqomBEJorM8or+WrDOwbogORpLvIFfzbNtRiKlgtUO4wqHxjQaEYRh15uQR7W
cixXR5ixFeqeOI4KdS8l9B3h8+oLV+5CFHyNBlCzGxQ5B13I9TEQ9gwu0eEdCR18FnPqVF2Ynad5
AXY3Oao/NV9tJU7+L9XPzfKxnoLm0gjIwOjRjcRZYTxwQeKcYGsbZRNx/Yebw5NXcUrD90QscznM
qFNtDImyBhXU0rXOsbs+YRZoS0cuaYe/GUByxR+vgLNaD+NzDiSuEFm6EfELtvtthepU365m+qaE
fY3/2DBViQwwTs6l/Yk6hPx3UdPNpI3/3v9Tusu9wwFzc0wptQw3K4USmTKVs9LLS+LsUBC0ikAo
nZcWoVWqRL3JNI//galPUcjxPN5jZFojhHfJy7yl9KYpLJ6ejaoJxkqWZxgYuz5Fh0Xouj1WbDmX
M9sMyb+RCRxjJA0lJLHXiiupDQGWvP5RqjfTBO1Db6tbD3E3APyxSX4VLZjIlM9cwpyafV7DRhJv
OKybjfABy+wtEe8R0KzAqtrhZAM57+7zsUoSDmUJ7lDZrcuNlmSzO/AIvwEsF5mhygYBZn6L5Sx5
UTSZwcD1pdZ4IMHXfxblgfnNYXNOEgs6zOYePyImtFL5euZlE9r+eQubb4pH9d+JwPFv1Zjn1rGx
25hIKhia9qQnld6m6pxdG8KIw31plVQcrmLF7gBCHRBInAbVcAjqfkBWG0y++SFUKtWYAGB4O54j
+cRkIXopCB6cas5aD3hJXtZ0r4oRd/e4SwUYpAXFZDylbat/pZVhxsp/4OYKlNj3N7CIXVw6Fp6a
9qY2jSPGJBvrXuzCj+BPmtNt7NaGhz6B0c/wo2p7owURq/zYlQnhP7NEYq2+k5tX2zVZ1ManXTpB
5fT4+IE/BzTY/x7kSLUwqxkDls9ZdzU1hMnLjjDcxIa5Qbp3AnZWtuduuoE/arghtDlOwPyYh/Z4
ANGsNPZuHmE7Yd4YiL35r9PGl6trCRJrxMu7HVQOLjh2B20GXhgzkNO+5Mq1ynQh0zKxhUocOlew
z1FZVUEjz7EJIZoDNoGw6vDd9X7Ls5hWt9X6u1WDGpYfEaCDPf3Cub5aIzjETBzffX/IDvpRKqYf
9k2/gmdLbfCeoYC8WZSHGkpC9iMRyHNGMc1tIUyjlw5dzk90BXsUY9tsWCMFlf66Rii2Hjsm/X3V
gu8xqdko7dcqekFCS7lZxMIh/QDM7mXueiJVUE87HdQFLkvPV12aLnjFoVPzia/ogU5OSFq2jR1M
UnQbFkhdqB4V4+vnhNRUs6qFGq6x1wsMGBABS/TXD03QcTsGdGQ9PKwT5Adq9T7UR8N6H9s9mklX
RUnKpyThIQofcCbwye4q5D3TwasbyiCXtFVOG2XDofN+Hpyv3dwXxemEwtQK2iwIrnPCyaVEnjBB
Pdi3UBMxryYd0g/tpOIFWWOOrZt3DQGUYi48Xo3AWMDMRQp1Q+x58AOit+WnwgrjDpnYpUfKsG+E
QrfQd3KONyM8s8Yrq/AJdpQcKhtOpVOiUmd5TAeYfYa60YR4E1YaCq2RBdFdJGKDb5yzH5+R+jqr
aHJ6DcEBLHFrwBA+QNQX3ad2rkXFQp30lZ4eRTX0bFE4lW1VlPvuAQcREC5OFHfqehg8La0C14bm
3RlOIn6PyQKv8zqc+NaxrqhssK+j/PYvKPp37Z/1iv9INveNn53GouGkKoQNNxd61kRmwDuKtO6Z
FdCoKxvUhbaV+r3fM8HoC7Xz49jya7EXlHG1xXncFW2/6BhXVQ2FsrND5Jqg7/dLF1yC9HDdw1qK
NlLSQY+W/flcrVyhlT9euwRUqmWix5nQCKlZUauTwDZFPK6D3W3Jii+USNkNMTR7Ic7vUh5lcgql
sXbRpxRD2v5rn/WWF5RXZgAAn3CgX0kkWfbpQ1Nb6vLF3Avhx0r9vSY1/EBelN2ngQ1Bc5Yn1gpA
TboScjwchGnGGONLZQyLEMdl0y+aOgLJ9MO5cRu1h8Kdrfqyxs6hEbMs3ORGaOi3pl0B7OD84wf9
/315BmcwxHcFHiX6rStknQfuLHBNhlV3/2ibDHuEEm0rIzxMSfQGYdzbIgutwarPOhK11pzDgyVc
QVbM+/Hkcs1sdfZvV6eBWXxvooYoClzVVpY6dzRcismDOd+Ggx5kgi157eTj/3H1ohy0ju6M0CFw
hZ8TovlbbsHA2yJGrADG59I02Phh1NcpV+YAlc+Jenv3Gh2Pb9/Pr+TUniF27vIOUwXH2JIL37sT
I0iJp7ry0j1AreATVuQFxzsBPBSqRXTGwJ6iKix5kQP87wWDcPN0D+mNlszAZIWgGNsxiyTcsH7u
/uImlEFp+rOq1PcaSnpCviNSz4kdXJjgYYxLplq/t7/Vn3NzO+vklL7rlTJXX6qrDE1KXtznrYWz
+3/m6lbzZDjfpG8wA5s8BB6NA6GrQKRQmpZVxPSYBKcb8k/Xb8z2OQKaVaDzEMsazLKvucps1jDm
55CF5MU4mglVSs7opXy7F1wVHt9Dr3giBHRTHHZ23YRrT3d0I9zDbcqNI1VJLniKlmG1K1ks8jfs
OAm303NIXrFHt2zo6UkYvi+tJF6hfulknpcwJ/XCM4f0WxJNlGGOoXB4j7aWazI5Tj+JNXj1QykA
WpbV+PTMXmKJtTWBY/h7Tf7LoggTGBOcDo1NV1Y/09GUK4nLlsmZhCk83rA+CfIN2aBArIHoCduJ
Hzrr3OosmbosibhzynQiPSnYvAh7DJScRE/pYSvCaPV3Lhn1OuWQavdp0QVSoEOIxif1TAADGgSe
FkH76haGK7X3mLcvrqgGengq8EJ+kWNfmx9hEjMUW0NqW/8Zg9rE8Vj1zF5xEA6gBZ4wvAxMFmDP
eK3THw5AYzJwMXD6A6V9reRaDJT6ojO7R/E+INmuveIm6vLtNTvLAoOJS1WP0KOZjHgoFDtgTA4c
I2vlRf4RSl4KHYU+jPiC3DetjkhbXg9KM+ZySE4Tuy0Sc7/MFPS7W1+NcwleofH3mOWyhYSlvuKi
dQtjouaox7E5vnwvKlu6WDmnIt53LzylSP8bf7ldhh3ZmqG7fXe5fMboh2l9sWdYOljj+W+GCSCG
63//ap/liD/SOu78w9qJFgnrQwYFjoqzv6kRJICWRyYLrdFb4fko6aP02CWvvCODmhB9PFgETSJF
n9ZLHrXsQb5pCtC6qVDbwSb3uhxPZDXOvqa3PrWzopo1DEXKfas0CPUJHSyBVpmUyF8AZjr1AWTj
KWz2JikIZlsz8RkeAFozaUbdiFSk1huCaQ4mzuV4n7mtKQw4NJsCyle/rDLhU6CVd1wwpaU/UwRc
N/8WxGejloDmA2VJJyccZHlGf//m0E4e43ubdLjHISVqc+TWC7nb0wAiqc4Txt29chxsORGlbrwW
HvaymE7M4Mt/H3LbM5atVvPBE7CDIF9opMQAtIBm9z59uh8drLIpqVvtl0Ua2UV/vu0B8N9XYukJ
haX5dVKobShkkQwHKK3GTJ20ghPEpO/cvhFQDMd69/snstp73cMWRmtgbeFX/92bm4IF9Ib+9ZLy
KDs1CAsPwgyp0YdFEfBWCJDuOIyMGtV7nImsIlJ4OuRRiXbgl8LqEe9aEg0JMOtUkyerlXTsgjpG
EMpQb45e3rRxQm/MH4r7bA4jBZCfyhaXNCb/c/lKl+G3WWkw2yHfbOpd/apgnMBmgAZFo6TUnUYj
qa2Q/kQOAU2nZXymRdE6seyn2rEHADOqAo1Eh37M+Ucqi5JnyEfAKiZOQkXE/kFm5mwv0p6phsLE
UdPQ5hQZjX2vJXmlXsZlc17VKDqT2iBTkrxENaXMwqw7IxTezjWlj1ZYxN1+MwmXxRrTdXhHVgVM
orgQ7mIJXc2XxWHClnFO2MZzlfHGs81xJiieM9yiHsOQgACWNVnp1FASf2dLbrMss3ve8EvFrBU2
zBIOubihxWSh8vZlFEBMBSOnn5Rb2XZbdq9UiedNepNgqPXV9+Ktv1WQ8mTY9/ISFqoKv4q8mcia
T0cx7S9EStqlGpLczSoYpTdq/txktyxl1YAzuUyn12VMXBZrwd61wAy+NcL8oW4yv6WUT0cDBjsv
lOnyWofjFeX/Mghk+3U3w5lpP50iG/od39fMiMD/aULbXJFJru9Zadiq2Ft5dovx1o/i0fnq/My3
T7NeGK3JCSEcwPzpf9sYiR8g6XtQGfTW0UoIyo11WNoICcJn20Zydzq4pT58TVNyWQsRCXPivxXW
obaGQErIAghY7aU4WTBvcxCc8mVRypr3aLtsvpQY12eepFluUcWXACvbog5mRGG5UalzXxY/XY6p
gtpnicWKxChWp+qANCesVa/QCBD0a7e3XQrQ9hUFXCrFABgej+wjp2v8jGBfC8qngRxvMAX2lVuZ
G+DgjwsCFspN+Edr2rIbwPdAgu3BjL52EmNZpsZOHrievB776SagELardMssVmboSnX3RGG2XRme
OeZFupokO7Y3DkVd8ORyw9TxXj8uzPw/VHHZ1Kz+AxeXBKXkcFBFSOTQsGQ4+6H7DlX7PiC4a/xv
dg1hK5daQc96iwAFmgFc1SZKYwRBkkAQWu4HutlZ4FsV+q+ShTQzJpcwx2QFLrw+D3SBfs5199ec
rl8ZcAaZavQaDdSmdwwl+uqFKeW38MQ0NTaj3fx4nEhQR1bd3xhRkF6EF4sFafbeKKjPaji9k4al
VlC+J1Z9fppuj5U+E2IPBcnjlM0bcvCWujgoxu5TfU9OW4LB/m7wyVdcrw147IzPH0fkCdmWFrav
zlmlPZi5cW9OvmzFJfAg2GPMyZ+YY8qQfvIYE5gOAgjRe6fPlC/tdJkP2t+4DSP1Sf4Io7WagxxZ
E7B3YVdpFed86Ek0PJgGYTr67knFVgRa5BjtE/5OEmbLUu4zAS6yu7SqrzStgeooOr32HPVjKi7E
h0bGYiHJW6Iwp/xZd1SvleTiEhqvFmgCaNN7Fs/oObaE+UE8w41MDTgpoT7s4ggyACFBn4fhSgFr
hqvJ8FDL8lI2ux3Y+hgUvS0pgpPywbkZie1KHXsVqE711rLit2dVjE6mHxZTxRNP4qG6yRKRYP8r
FsVdvp2Ax1yG1rhm376a1id6wlkly1EEZFx+PxDKkUuIts6eY1eHMauy5pHXMq+3SqEgNURnq31N
SxL+A0BaghD5/zOLikeNYpGxX6NytP0GD6M08fRxg+86Xi9sfBtlOq/Atr3yCmZcLas+CBfHSJML
8jKPheHIw3Nm65TjHboSdwH0djkbadGZ0cCv3bG/adR+iOwdjdy5Q1ofP2lH8cYgZr6dO1DB19eC
OZl+H15hwuCTph9dtEsuSZG9+PsJCzlbevFBaveZyqiGM15NnOP5E0GzJit8+PL9Y1JmfLfh9PxM
x41cLTxO//Z+Q6cSSF9bmBrDRv/wVOfjzxqvXjfYThwbzB3YNsm5ONegg4iG9FzmLG+MXsq3N2Bl
tSEH2R9zj+p30cHqORNa+ssfFhJbsAsrqhFKJ77p6a8FarBBGu3NhYEd/ulMlB548PsJJhbzoKfN
Ngh6X+vEcxMXvspHUCE7QwIX/eYWyhOqLJbWt0M73aZH+VnWCMzlGB0AC0ygKA67g9JuLZBWog65
jxWdrhBMk/Kv7fGas+JH27IgDY9S/3dWF02kbvN31ZKurZ7PxRyw0hKk8YswU9nh4m2Q6et8g5VX
492lDc9oGq4yomYR7FOSXGazdHErhrmM1Fumg3l334JyZK97rb/2ewbFqIb+PbCXRfIU8FRWXqTy
AnyQb17vz0CGCLPcaWzTGbqAEGLpbTaluqUIgtZc/4t1E2sb11VpikKV+9ufUodgHzBgqpnCHO/9
c7graKlyV9POBZlHe4Qy2nkZ9e2cqh9IXXNoC9UtKWNimyCQaY0Ajy0MpZwVboGf3DlVFcm6dWld
QwTy9Ai2AoNMWoentqtilb3MTDEEjRbRVLfRy38G1LWVObxh1AmImeKE6A1D5j1Tdd89gipoXKTK
HdQ5nLjeTMkWksxOpgXWPN7AbpMrZWxGX62SjmFWQ+NJTlao6zZS9udKnVo+NFDHZlaDByLScE1j
J3YnHdqiqZ41+ljdxk/Cu0zljHbKcRYvtnuefffi8cgagu8Av/GwM3OBgzGjVC2U5BYA/vWMPwXU
6BV90s28WCNkTad2blSCIzAga/KybLzK0mXTdFKzkC5gesi7h8bqyHP5e1FBDCt7fHCREYPbdv4I
3NgTCQ0ykoaryxzK6dwhpWVpuCzBwQRXYbzPlXCH1uTnwWHxSEp/rUzK4YRBVAxltzNjudEsHX2b
RWeNXARz+ihtCamvarZp4iDu6EYDi6hxX6dv0Nulxf22LnUA2IRDHn6DzIEjTRIeOQWWqc0Bd8jJ
IIC7ZKIIPZ0jYkQkWOXJAW1oI5wqwQKmCx0KTkDff+D5vP2WjsABwxHmjeGh2+FxLs82LWHSpocR
IaxXiHn0AiftwgG0kE1naBNuvvqpUib1fclwjzKTrXnEItSqUbARUdkEQQgTKJSTT5uqj3r8Uz6F
SZssCmG/yLjdwKEaufbqab1FlH+MP3nvdoiRAm5OovgxXIr1Kh9VrKvqlBaWWO27J/a41W4LvWCR
D20xOhu3K3SMW9g5rnnGNd1ClZHi2XNQs05SC2+RKvhG5MiGGfH3mi/zycc3Y+Vtnw92dEcmW1DK
eUU3SRTET3sSvrIOuD9XoLTJ9ceDHvtuT1hXkdiaXCiKNkwoTSYVzq/3hHIFlsBcl4a4VhD6qdmx
JAYw3gO3MhSv5QsZc4GTBR/isN34cc1Uose9LSsenGnoB+R9IXzxRz2POB7DmYU+VsN+bnz4MP+C
QPD0DbeAR7JQ+JdqFXRcB1XNhMVx+P95vAomkSIET5rIHJUx8ZccTPAOdqesTUD6niPQTZCv8/Xa
QEZbdsnra0NGeT5wxnJ1wBHMsB2etrvkl2Nqvu7ndgjXvfW2mp69y5fShYz/zg3ofCDnCP/dsCP0
u+u5S52H9Z3Bvi+5mpjSWM0Gcfky3/IOlEQQsSrScvwaI48lFOeBNyMYlEPKpnhohgIDxdGIruom
YDNXk6dCzeAd24c9KtP2C9DLfhDgcJiIdL4uqOhgiV4suqWp3Zup9FV2qrC9Wc4Ke3jYIHzmdCfu
aIiuoi1S0HB1c26CRNLQZ/02GLkBp83Ity92oD8hw4LD95ZCx89+KFmFqx2dmZ1f44i6vQB3qkcj
AvkdBMN6UhAWySXE2wSupLhaiOtqhdS/K57oWvz37mP9DnlAUdrFoRZIxNmxdDcjaN61/95riUJo
p0YI8NlKjdRQ85zJocw9pOpJ3ba72WdkukXJGZ10cYvM+DmII4EHLJV7cmTfbhn/zI7SyiEmoF6k
IqLVN8g4U0sH0CjMFBHQb/T2hhMWV5kYkS8CWLIwYfBmvC7BpdWKeO2vqIhVQsr8QzhMV+NQk526
eyyD9jK8avHl9GiuG9gSlKGXw1/690lKi9SluKcArGjrECBC+/GHKiEav5Y/LKNYKYRObY89plml
4Z2nGlxAUWfm8AMXIl1gdpTvAE5S7gdpgXHmDE7nCRgla1iY7Tb5dDjXbD8HqR/wEeh/XEstPKaN
W5zww3v+ANEhud8+6XwQI7yKsyb+CMVacWo4vRjlC0PVc46DL9XPzOFhlQ5m++8VX88FRyUCeX6N
DxWhvvipuz1BSw/b/6Og3+cPbCCWi+dtxr1BRM/eQ4f2kFTPqSUeBUyCDulpcDaZ41wTtLW7/9NP
vvXVPaoVtd9iPLIzPMXUdp2Xo/vEVvuKQs74nVQ7A77BBZ/m0XtP1bV9kX/CnEmfvYH8NoTFOX7I
u0VNOMQK49hnA73TqcN6iQGRyBd7FQU6job0QJWWyvIYoFg3iNgZM6LJCj1KJujdhF4Jdv/pAVfh
cWJU/5FxnDbEiWWFK3IM505boawv8Q7vYydG25VUEAFuCWPqOopwX1PLgRepNzRIHmXLEDftwOQ4
g0fEMX/N0/9c/LeNfNXBzUHLvvcIdWiMXIcScNR9oj0tJjZ3aRC7hPd1QXcWwDWaeyFJhu+W4I9+
WevrsEmZffAaKB49EAciuVTBiSqJivjz1dRAy+SZozPd5AczQxvY3ZvrS5gqt7uA+LILjKympXNn
ssgKmAzOWLYBATTd0Qq+C803kmJiVH3D0YXG8/Oa1Bqgj0g1EA2EbIl19UeHeLxQuBJeipxVoF5n
/C/wSCBNtZ4DvohJlh/gpQIDhbaJJwIvmx6YNC5ChBSy4a6g7QG/xFxWisswVkgnG10CqKiITj6q
ozSwxdx0JLO8Oa2HQh6GMF0vBox8OkO8sw3d2gPdxpXuHrdOUsyFNPCOJwzNPOqkVgL5cJlHOLPc
A3qFNtWuwzBaYYwkoqjIFx7JLyDkNCen8rpbVz1JHfWCYNJZbyGOnoXrERM2rpS3Juq/InDXToME
8CrnYZgG+CQqsCKAaK8agWv6UmHiCXsHwzNZZ1MjGG1roGZUSDYzNxN48U2w8Se0CPfxu965ZAbO
ETkGQnFiBv8cneBlKKi9yrzsYJGfUAVDJjadafuW4kJWM4bAzjq2SvtaskGZ/uqFNTuHACsQNtMg
5ayO5QKWpUR3+YgtN7yk09Z59Mz7N5ktdv0CP0Ij3fcD5PAS5R3+DmM7BuVZygma/LNfkc4dAfj7
0UHVpJQz7A9vDerHgsQaOJRPV331dOW+bCoaoQD8RqO2Sa+jZpRkKwwQdzQu7GMS8gQBdYaQ9ir7
VQqZ1oyk9wufWO3vueRgHmkV5VtFTPyIp6oDjsnxZs3swzUMq1ZlUNPJgKhY0bTeQ+IXUQLU3czJ
f5uLPV3aNRb543xurr843ydWmt5aXlKX9/NSvu+aLLfmxEir+Set+4I9eHVW+brwXoPvkNZ4J2YK
sC5eGvgUV79lWjWz6LglBnncJWq+KqwLvWzklqkDgy1q1jObx9rEhOjwEwV72mnrWGr2OWjcpxG/
6hxDIXTbGRH17QS7tNVykjnLWHNKMqo0zUdYmw8rreVw1Bks/Egch/smUVg3mOEwCJKGuGpFU0WU
WuQUnDREQJnX0Kbn7uQcFda71HLOQoi0v2H3RWzOKuNhATPU98TI6IGzOuSxfQ6U0KSJoXKq0xpS
4oXxOM6mit2KClagOgd48/cHfCfzPlO1N2IQXeMOKdzC3Ie3S2MmQ/87gLEdT/U/2/gmmnhuAz5c
3i0TKgiLYfHzR8V+Zzml0O86m6niVrzUYYH7mXoj2Qz4/hu+GIrBUeLaj8MCbyXC9J4P/q9aOJuL
5koTI/qWK8G0O6KIv6aykRJGOx8qP1ZOvXi8tSD/HUd37ARD8VWhS8gMKD4RozXe6JVlkOuCP0ZZ
HvB3an2b9NS5ZCQlNIvppeQRH/vtwr8DPeQzNm4xIWk8B4a1XtuIHjAjtOiE8j2JbUGgubmfp+BO
okbCqefMFjPFI0mkH1UFbaZp8Wwuj0neDsQqaXCSbszeKMDJIXJYv7sJ2pcokbFMsGKDDjuQ6fgN
r+tlna/sX3xVb/w99hgclOFFtAHXhOk9kbR5tvCnJJ+TaD9S+fstYgIurymN9kcGYI8LT+lZ5dSy
0q+jsp/8dzSEny1YnDDnDda4SlvUpOXSSeJoPgMhl5sPSoHHidxHI2+WkXWR4gFF3RhtY4ly8b3C
0W6YJoAnNrvjBKkJDF7SxrMQ1QHMV8YHZSkeJxtsr83qneHWzLkpqXLQhEmiBA3nAWPRazaGlfL1
4MYwty4wwZ+8XGOp9Ihp/Gmgu/kuY0XVmTE6YUSkcfmwFSm6SxttJjcDR1Q20KhUEOQyJH0hUucQ
SGlP87Asu52EkDjjMmA9SZoSjMMB7R/QJboA5QtMS8Tru3Aqus5hhdFoNh3Ha+N67WwfgCyEKpm9
Fw45Z8gMmXyRCyxJX161pQNFXVTX1kTRxosPEWPW56yNqN2pHjy6WtL6axKNL8GBdpv+ffsOjTG2
9mJjF3M7kuixXi8e7T91xDZSeeGp7nFjJD3lqWylc4dSfXZtNfznZm43iXtnocs0JmkWEnngfI4C
RPNiZcTdGJ3lzU9isOjPvrcU3FTLd0mbaj9qNFwYWJLIpcIV0sudRBdHVYuU9R8aJsM4uxOMhyn7
6sj2J1+Kt9G9gSUsqgErkBti4t1lqQcy+LznZ2/A934Sh16iyAmMUiy6nsyvpxgeZ5pMLmmwt3Bk
GJOyV25UP34n+PIKzJptZNZ2u5GxpxoVZAHXkij4Y0RCw0ZzRSRDEMcvXgH4jGb8IDnM+mmawr4b
w4R9Ter6fRc28I2BwSegiExb99ruuR8n0PmxOpYG6Akz1tZSxAIf80ERLG9bLN+7JiY+SOxp8YDS
71Zt6Imhqmlyah72BF0B+6lxbEm5RrOUaxKavbfhOJC3JSIPju1I60pXNskzqL+l/9Vc6oL9jlRL
Fb580BJIquacMNdFBLe1XL5TYvcvDRbusH0wj2VFEzPBqVTQXQkhAbHgdMu5Zrgp9yHZaRpKJ9sj
GVvFDh/ah/qXG1B+ZUjXn4v2M3QlQ0GuyrwUnJPA9J2tf5AdSP5jogJrKrYVUMlXhOlZKj+BG3Un
q231fKhhdCJwW9hMrP0j945OievforSJ9qYhOxIzBt6skMdp2cXzsAs0wwCaeag0+LMawD5x1wBi
AhqaFt789w5SEVpn/63+sY/BaAKs6x/qBkxi14ZpD4RJ5zB4XfLrbjOwSi31jafUg4g0xGT3cHBV
kKHy5yrlIoWpYpQpIg7ZiB4xZHhywjv4PI6Eyj8MKFpybRyjbPlm2eE3U9r1Comkh5wlHyUXCf7G
t/tYNSlCtkIrJP31kII7DaatKPQftiGhZtgNkk/VJQbby2I8eHuc4pIu6bbvz6VmLX2z8c1nB7rT
wTiWBpV/+PfAnr5iRfSy7a9YVBxzQPMK0+gEU7SuPWJkpSRbZ0cOwLekE6wixyZaVqviNoGNTDjT
aSawufHYeOoBmZQC701a9+RC9LEvcv7rhWjBPO/tCS0FdwknY7q0trttWeblGgtp+Uy9AEbNndQK
7e93OpoJ0jhoRqWvw3VW87G8vET3WUpPGQd6zXzSrNzFdqDLNm4jwdTFNJZ/iGhQsbcitRP3+vJ6
t0Sw1NkTvgHJa/KemDE+HkFlXOv1NkQ2k39yBXRg8inXJhJ3z5JlXiyRqDxFMo4ntYMqN7RoQ7Jm
bMuTNBy9R6zvtIbANL/mZqpmvz8qISx8JK3EawVdtpsjK8gTX6w4a4XAwqTreq6K8Wg1ZGCRORpe
124g3rK5oc1FMtax6dParXYvWYBLPvpGdYiUorZFcE2Vmjq57cFTC69+UpMP19p4oNEnxjDrtj+r
sqHO7rJ9JsQsNesSxL7kwHw/kpJu9AvYe29SgAgT74sTuk3rEcpfJVJ6dG1KYsMPJVy75dfyDEzJ
iA/D2P4LTseRqZFz4UKC2zOvD7V84hiPVhsb1V9biwcTDw94x5XXFzBLC2gG0kxWWhXbIfWQJWMV
SSL/ODqVy6UKgEBS+waaKKoWLOT6t6AXgBQiW5t1+Mn6zK9ye3GccTkkYtclAJgHs0NuA6CMSkwG
TGqext56FMix3YVGxz9LorjeKD2Cfey8SXLVuTu4XvBvssRc2ReiUuxSARA91X328R7qPVoiORqr
M8iArF06Nx246X3P+WSdFAaqxV7zYIP7NOMUi6pWME40vsLz7isVPotc5cqhGmxQe0Unz99qn5jZ
fkeQcg04vgxK2uYXRkcIrg8kls6tdZ6KNfNJfUDyyv0SwAX9fe/NU+bBKFqQQ+T9z4Hb+x2w/2Qh
bbwgTy8TMYvwCE5pgKS4Hi50ocXfkmoamkg5baIbtO0qUZuHwThQ5btoLN8Ho4cUTnzfS5yEJrpo
IsiV0VE7Eifqb6i96too31sUrnT3AbXY9NzuFKcD+vD7NdMkBn0eLyD/uEvYmbiXh8i5/IW6DYVu
2AeZQca88w9tGcgUK8gBPUFb81OA9POuPKxJKdesxTtdKqVFOwu51+648PVpiUMaCqfabYjiBdpI
FAJ4NNkyJHIJHDTIfurroh/24lMI920pQlVMmlf1k1uMGjHRiEwhcl2JJrNCg/ZSQbmnkbRexRQu
vWR9ucm6pqGDWQZn52mbp/HPUzL/2ilZ0fA79o+P4ey+Pc5aPSrzmd5yZzDoH1piSljUJWacWzS+
5e61W0eLprM1JivF0v6pZiMypoz+2X63Q7x2o37RujyOGjzsz1h6Y+CVHH9Q40BPE7cS42PSgBHN
JfpPRZRWGtWmeQGHVMGQvXRlUFVj2xE4NzKPFofMCYNv+SWxFqCLZp5XHjATYDxaa7CEvgFwZZBp
16tZyoXO4fS9erLRdIUHOhL2ev4N8uybNtHzrSXpL4j0m4xi97vsTfN24C2go8xHJpW1jdjnunn7
XVZ7H1tbY6+CWQYSIA3LyFf9jAvZYwb77j8AZI1RSv5hXTi2jhES6EKkY5uwSH/vyK/v37rFUPfC
q37Ne1zP4YXtT3iWUkNal9W+m/98c5r1hInqmslllZS694vJM8APxk7E9Lf6BQxMfhZCpIJRrMkg
im27P/YlJVXdDYJTQNU3pgXuzhjAo4s5iOwc8JP1ggQGl+Bri3btwA/dldnyOEarpNBAv55rI6Xn
eH4kRZ5PS+t6wIHJ0C5vMRxqVPXuvuPCwykS0IlFPoiv7jcb8ZC938w675z/QdES/GfM+es6rmBW
XnkCh2C2kpNxM25XOttQM5cthzxGwQcHLBm913fHJ4f7adfSukNS6gGIyKRXm/ysImrV5a1YDGYV
B42P4qLhUEmtxB8eI+o7rJ/F74a2GYlIxym8rpT26wIvQnCX8xcjUEiiOm7VDpXz4TN8fuXC+h8Z
VtIR9G9sRb9X79AuG+26Q+z41u7NbFAo40OVsgAdpufdG4rGbQ6ZDVyM/Cszj18SjAjiGsxHKSoa
MJXti2H0BR20r4HQnoXP4o+Je8JCHxCPhyvEzdeCWhist/1w28pUSNTCF7zVc1krfD+UeApBitub
2EMoiLe0uuoJBQkseM1UINnaqs5QLPfqlVR1zrgKNxxO7HWbW3Ok9oG6r1bIqIenuQRAewV4YtgU
fnJ8ETXIAw3IhqkGrXzUocAwhJ1/wvILfdg1zMSDGk2rHR5MF8vwtFLZmNSPDMYQ+HwXgJC/ZGOO
BMllgGOKMO3FqpC4wX7ojRtfgGDamAIN6xtSCZh3YQISnBUKsx28Xb0i0R96yJAYC3rGd8/S3jlc
46LdJmsMqgmqlglMQugXLYqeHa5ta7PIKrfIbfr3eDCnVj4N2Ix7D7dfP5GrklRkV5ks+kmgqmDa
4+8BnQ6FCXIFCivBiUEzKFYT3fzEscvN3Oe6NzaH1loFE0Hvyi71A/smfPVoQxHUllurAUb1V0P/
YJhdDFqeh+Ar4Xvo21Yy18SjY7wVzHv+VvjOUlwblLg8E7HPJprl81V6X6u+FQH7TPCPjDb7PIkm
C9CGMSl2bIuqt/1GZSAXkjP8zBrfWH7i4XePt/phzruhNMj+aDiLWjYmy+V+3uUiHD8FJkW4rT1A
jYkD6HMFphDwFhgnHecxnCOuYFNxhXb/dWuB/MSDRpn5W7v0C6YhJS1+R+pkrssJYOKr/DRaYM11
F1KHn0ba9EZs4vVr+9arJVYpe6enIHX+y95bBXqw4hyzifkNH2LBx8Phq/rdBULGi39WtXR65BPc
UwvbimDPVd2tYwLifaCl9oEdqbvlKJGZ6aQRoAr6rozzAGuOso5OwA6Nlao6bXgBbLUi4hmhZcG8
Q7vPGeURUc5tcw6UpUQzkQUA07NQfpUFUZ7eAeB1Heqo2o+Xzj1fMqhS5RefAQLg9eWDHif9Bnq8
iCoGCIl4iF4rwyZrKYA3Vw+IypxMB0yRGJFxThI5PqDSuTaQeXvKH4vQMwcbcQeQFV7/wOP81XRP
V2Yqxncm3iMqvgmLsWFuWDaiH62zZG7ooscj/jEz7vWnNInTfMS7wFrtfuoj1mBhHnfs5pRLh8my
wOT6V+MvDdTQfMgtO2KY8YNsdrkDxANOBqV8+1KhzQLfirv7mGXvx767IeG54QjDmNtC06uD1rqy
d/KCSoTgLrJpeJSNs66qdiHjHE6qTn/m5u8cL8qixBIhIcJE/b4Pz9CTZsZDqcfgc2q3q3zFxw+8
VfrmJyDZctq2hbdLpUBV5sT//uq1tsTFaz/LZTZtKN7NYMspJDTBGETh/K8pneiEtiQ1doBtxelu
VMWN97oMaRwhe3Y6ccweheX/m+fEKXD/+6Y15tQobyP6ItnFuxlIIPHtq9TdZDbquB3Nw1I1wgAN
HxQnQNQtqpZ7vFwysdOPxMShS9iyfYg8pnNyLriSr4budIVJm5BhSIYJpz22PD3jIqiKI0TpaC2t
FGmxQFLffaP3Vyk80W1SdWl+O1d/P5Ijg66sLFIa4AkFGNAOZ5/705ZLDdoI0c57FQsjIym3htHq
7ajwNZGAatj7NWfbjt0k5k/7rQ4niKAeBuol7wB+tHozYTV2VHUrA6RXAy0Q2AOrC0wjEXHE9U+F
7PKOhLI/5APbQUYD/BgFVfamw6wU3Ldez7VwhcRD6ohAy2V3DM3fD3kAsxZ+Ebs3LYwH+Jy+3zRI
DN0DNEV3YJmTXilva6VwLTa3vtjPy3AsUePI2WWLCrOxVpBtzjRKgQNrdBPwa2jDJBj59XQsB/PN
40Y//10RfjBE0d/FZCbQ7JhO107VbFnI52pZvF0kHHTjEuQkPZhcakUul0X0yKmoZh9Ufn2h60Ut
7OPmHIkGVSi+Lkopnf0I5ysDXyMYoy3gc5gtilTo5JiQaR2DiTjIWe4O98Swt8YXu+IC8UJu5Bzi
mH9+EUNYacFiTb77+A2uuzVWyLX553HVgrhoTNAyJf6e7U+sePCrr+4dSeTDnXoTUx/S/BDqkl+A
D7wiZshYpuW+m5iN7VkZkU9lLyzDrGykyT5KYS6/A7MwZBEl6q68uLTws+qFqKEh/AikwPeKt87X
njS5J7W48rDtyFprymzGyv6uo9uW6OY0iQmTAhW2iTxeKi4XeBerOJU6/6mg6oZrVB52OxieSxIT
ifX3+n2J2JD6fGcQE8BFnLzyJzEhHQ/KS1SaNKE/XJeppYAb63Pl9M5pVJ9qMrstQR4i+0YMlIny
hPzzoRwA1PF2eDGCOxrC/o865Pi4bRanNXJQ0eFvIDAMvdTgYgUMKtHEPp/LWdFU+v3S6um14PfG
cMwwxsx+72zCF8sH+ZkXvSUc8RDodAbqgT4NchP1a0UhPKMcoEq26NnvuJ7H8UA7IUBTrEl/7eQf
qhvdIJJL2uzlVx03tUoYHCIUdOgM37GM6N9+BXK7LXROzi1I1LXIHzR3EuwUH+RvAHOX4DS23qe5
fPBXS0DjKCdguZrgBs7PwBDcZtcGos1/l0Did3HjnreTflV6yBnExzrguL0PiYO+nKlWxGM+ZJwX
9tqCmWBJz33wfzHYSR9RODmmuMMXXUUknKialDCFdoQ8pTTLnwkw7AiWKYfwHe/2oerrG44HGuGy
xClqhAZsLbPFbUpEZ19Z1Ouzfzq5zm2f5L9+j2EhKX5oxStbIKEtbs7hJCufMSM7eWmX9y8VFXCZ
YYSxjOkqpEeaKIZY67QtPdPRf74fN1xAqXkKCPnHFYZKlPMTkZRg0PX7gFGqN5Wr3sBv6kMduwcR
n92ZK7kuXJDZA516NTBpLL8qHfpVM/xYrWWnzXbTFB3T/C2vVKOkmaKjRqJo3XRM2vnCBHu3mRhM
3PiyjBdcBZ59lJdlNC1Qm7FWvdCzOB6p7C0Xr6m7nAmCHnaPfULma08nCYsyPL1cDXzu2oEbbV56
cxfWJjWrVv7ap+yRaGrfuWKpvtKnAqZLvHvxRN494KyvUdaBA4tZUWJpjz8KpgUET4TpjjeJf6ai
ZIUcgpQGkOD7b7BZhrakC2PJkEJ8a9fT1Wvc5UQrKFCvJY3Z5MC3nLfxR/5Hgox8CC7U2OpgMaKp
m2O2dEobiGcQXfTGrC37QPOuN1GIQYKjpYpHQB31xgbXFKtEIH8t6eLsQhYtnPE0wVFLqpksWnBg
PIhMxXgWU+iewj6RVYnWZxnp1ZQxxGftrtR6KsEinJkbIWrLrJea+KZ0cQE4dhzsIjUA7MwtF+7E
x3FRQnIPjPRpeBXeLGZkNN/tVtokrJr0UNbIt+I3euZS7hslx6KnCDTMr4oKfnqaeBb+lUGsJ1g6
OKmwLGSIXU2aU5PRsDFEgFgP8IQZBjJzrd4FVGMLI5fpuzMRaz4tlxiM3iIpF/g086ACvvvHPPeC
WmnqnXtUyfhSUZncECuNL3HTnpjNpk3huiAoH80Dq8GHWHgo0lAFVqqp+GIa9KUitik/HiS5Qd2S
n7KGXXhhpQHZo5l3Rw/ddeCuyvzBde8eKSnh1aBWCeEVlEiq8iH8sg091xc7nW41DHH0C+3F7QtY
HL1WLmJ1H48km1h3p+gL6MiTKFIz2QYrjHEk2y24yeEc3B3ExI1D6/H7tN6j/+3iV6P3ifckcb/n
d2TsgRjvXJwugBRHvKDM4zKb3PXOEuw5OEx+PnFUSZ2S34GifOYHl8zAAP8+CN2tzbfCB50NTLpv
4PacTAJb2Wv3qjLMiytViUZUz1RfGlQTie/U+q5B5q/BkxF8g2qigm43UnfCvSls0EskNeBSGUlR
z7I584PZQeUxYRvOHDRl1xPbVKfyNUszEbH9NsaDUHg0I+sT7/Qz7q0Hy7zj8kJ3lFPeGAFMJVAr
4fhe/r5h2ZD2pxI7IvPBEFP/Gjul00YXsKrYtUEJ49JBZJc0g1Eulb8lXAoGfk5tCf7gEmM8jvkD
jIRr++VBg+KxWBX4/CEL39dWtTJ9w0dcbk273bqpxE9z9yMV/yH9lQaay/vABGpk3wvvC7O1N/0Z
FW6Qu2CD5bqrBCHfFvjsuX40rRbH/j6IkBxKAvepjwlyfWKoVssDGaFs9Hh4erVBQQuQYkQo6Bku
XBdL7lYcd6YBerkXdKSBpGVD29QPrhuQIVmczIq/zDdcpGruWp4csDgeiZ6jRHP02TsYm3qn0jA9
tR/iORzqSzO/4yYAdtkZ2F8nUZu5reK7WQmTTvTsJX5XpOW6dvghcIuJzm2iAA6PuKFeGaIUXnCw
oynDdmVXt1p59kjRPjO7AC5wWX+1lo/6hiZvtY8vxur1ebBxdqfuTOHKKCa6/OasiztSvjYXEQnP
BKwQAzdXIbE8OltwdPYhQa37EGpLqW9LZQbOdst/uFnmGAOM8kUGiGlGMHTqyYqXOXhhmCpq6zQy
xVLcXnCBJUvcbRew56KozJrMqXwr6AcYAhMP2RLnXcci/3BJGxFznrJUQO3TVRy60MTZ/uLiKMoU
zcU0bcleG9Y6jqtY6FmcBMwS0nGfpL5jtKVTuPGpXO8NvMvwzIKcmDCYoVVEt/v+8BNMr3ke9753
wA+Wq0ZCpvwA2Hb6Uob2CO5zmqzXX68Du6jBjouz/tWGmyI4VKCqcbh5U3dd+pzFrAZDJ9I6K875
5ZYNJHmzgvn04Zi9yumHmaGPFFzicZjSl5vH4m6pesjRT7YPHBLdrgHmMaZIexMkGNklrTIEHEEW
9r6MVj5W5/D4KlTYENUIRsig2JY1GJXnpqFrxRd/2J1FKbSK2Qqrv/aqe4GnILpYzRlTSLSyIKwU
WhxNxbIYzOqh90GwNAFaVI32f23xquU9kkD7zMZyF0IVwTuYXgKv4/cLlQYxkIajEaZDdJ6bLal4
HYkmZi2aHrFTcGXfbVb2uNvjoXRz4KLmFsyEQUgG0TIFr3eHMP5hcKKd9JGIeEScLBOeHbWAFH9K
uc1EMVUYWIaJFS3euHHsq1HiTV5t1Qln25msdEAFO/ks5DwUMH9eIfs+cD6fXZ28tpMTapUJT/pB
Gwi3koBHx0FcL0vkI6PNBX5nSBNCC1jpQXvZqEqIkRo48IYiK9N446Z9ZS+6MNlDD+wMS6saK2Qj
+iQsCybPW+dvtLOJlnAsVDyCRkQ6v+tFwzRQTJ1/Mqf54+hpsafvLJPFGXyEenCw3JjZcDBeSi9O
a1LJVJHdgRE4QbYZXJW9sLJir4w2QsPt7cDcbtiqNMulAoyM+RBQlsvcVgYR88Ob38UpvBJIrQ1y
JzWcjnkVogrxJihpy9dNh7/gmrFx6+7D7o3pj3/vsYDT8vlU9cgK2HfSS3yXJrYQHw8CXeGO32aC
qT8bPdz39wO2zhmTdaFhC31fZywxt56BCD8DJoU0MpH6wIm/SqeYgZKiUhuIHeIm/ub+r2auY+FL
Pg3mBbWmaNUycPngwqLjOHv7AsRtP3fYL1mZx7EO9ajd2tq0wRrCvPmg7ULgnnJOjOjyxSgrqpUY
rcurlGU5Y1zIlzzrNNH+BGiFpEm1Opd4f5LeWjBxnP1uLmfExCNVMLo1FhoPif/+Eh319ganT+NY
ZUx0q3eA0GKrDfdZMn7C3yi3RJuXQh2qonCnPUduqpRVaEZRBWhG9nOa6GVx27f/WpgdsJzXPwiH
BknI1Bb++PHKo7p4iOjc3CWVlc//7VRxA2FqozbGjuX+b/oqNDNfvwljNQ/2knd0JGXW95cLkMi4
gJKppC1OGiml184cDt/OR9/abcOasoUtqdeU5VoqIFCmO3fvZtjrTZz8kyyg6nSBY73sqyATSO2B
O4iLfya4Xx07fPD13WySjGMfeeEW8uEu7KtdjyLBJa2SIpLQgSdFXKjz+vY3FbD6xw4zN8xg58u7
xpQvuXepj0o9n2Li+Qlf6M8sj4ooul/asBE72YEg5nzCVABKmTnz0CpsAJX6Vm6Eq9NXuen3ANh1
yWpSjd8YkWZtvllAZtXiErkmL6OqC7IFznSfTVayDZyX/T6WmMrCC4DpW8KM/To8ZGhzx6pswfgq
v8jfY29fry5VaYheMnqftBYvjljfSz5+lZwpfjjrvnaadgtugmkbwLc+Aqu/8hucoSj/fZbBkVf6
pU8VcgofWm1JdUE3GifWHxPy5tVGdBQvkaY3P3eoB99ow0MFDsP+OBa4InrP6qmgpfOgvSZ4l57e
AZ2hay5sfQrwwyE4H2RkAzsh4CUxQuDofSpL7mfnWLBU/YPu26iCdRNywVjfeTdCQH+ggJjUBhox
g1V3ybrA2dfAo9WxxyHqgemWr1+ivp6yFSBx/HUoSYy9oOafAwJ0i8sYRE++9i+8Z8FZvWpPzaSf
sixwzTz4wXygDf+0FUK1RMf8EjccAOSTyjjjR+oiK96dIFGtsnjC4tN6Fx9mI4x8hh1fwl8apC3r
QgrJlD2fzgfu74dewPZDySjJksbduacTYHeqve9afVuSwiCEfOW7Gs2o6366EWAtJ4nAfsWBVheS
rav2jbrhoGeRP1XAufVkDjWnhfdbAdryFyMy6N3BXZYxe24HUeYVugndHThE3irMoFUogFLVIPvT
Uzv98at7FAZ05OiYvBjuLBpi33tR+Q/BlT6LQes3Djl/yU9961tr3IsFytsDSn/u0ojeueOoZ0sq
iWXYfhKEFCC8J6nh6B1P4tDwerVe0m43bYLMLxtsfqofdKtKGo2p2JwmxuB9cn6wUwvHG7X3Mivf
F+8DpLhUu3+LmbjOtf5APXhspKJA55LJ0qSTwRqD+0jLheL4P0UWphMCMevZdQEx3f1DLbly3jOn
8YC1cp4aUz/3mNRFW3Qan1in0n6pq1Sl9YQNz83PHitFAVTjdtYUHsnl5FlQdr6BHOFQNhz8rrKg
C8FdpP1dQxI9eNyQ35BOHanyQTVJRikn1klSpfm0QVl6DZbsSIe8kT1REc5Gmz9UopQz2KIhD0QW
NIRsneDHyqhUfsAwf/Lr/ftIwgIRgxgUVZWDYm8eBqeJqNN0sxFrxeDoUajdeyXxx4c7UgVFNg71
EXoTqF0bq/EH9UAjJwW2Lg0cKXnZJXTF2i3h5xv5QMaYNiQ9TWjTdTt8Lfc1XJqjyTNxUsJeIZ7q
/SpmVuiTYHTixcqn9qwx4G4j2vxEYFto7SfnL9NQNVoAacKGNRT1Q2x+r4LSjZAmyY6H0EH80fxo
0sjAEZIXidRb6/BLOO1r7ISeVttsJGtDJ2jyR+FYfBdtioLBIX0WYtD+WYHGoI1Q8COJFkG8s43l
tPnX+BoWB/15y8f0cVF9SRWga1Xy5bYIAmNMCRRnzaeC9e5VdywLFs3QUVhm4iAJbPvlCEClpZPG
TShGFSGLRIUgjOiQw+/SuZHcwE12TSmdTC/pGDrjHAJESYxH00ibn3vq3ZK2kJLs0PUoJmCKY2sp
CVwNvET0awSPVK7OryBqp8b2ltLRNjtYHmP42qeOqEuhkksMt4etuCLfIaNbfpjxyeEHaNfNzIvG
JOswpoI9GJzMqVrRAVOTHKREvFBUBa+m3YV8Av0xraZcXROPYOFrg6s9C2RFyb3WBeIZ2Du48XZz
uIjxQbC3XOtNmte9iO2LMxz+SwghKQPHoZQWp5+MxYRnP4oBnRsJNPr7Y1rag+R6eIoWWBIEUsXM
wBCrSay53lEMmHBfD98a/PBjX6vJ3JW1kBxg47XQ5bZ5sGGOfyQlRlF4LEX4YfiYJtKAVwWZ0EAh
GQGCzAKzHX2JUKuLa0yLRtPA9qgZcnMO3odb7EOV/2Uv/GzKFXz/TQfFKu93SkPcdjkpsYy/nDb6
uMFF/8bzueNcBDkPGprZyrdcZpAhjj3Ek9145NCQUIiv926yGyAPkZLX10w1Y60+3amad/4PQ+LU
j3TiKnfQrdHOnExxuay518uPCqWZPAXeNbjKi0xI1WIaMI2PTAAnEH27HXTkCfo63GaA9vMn6YZd
5U8froFVkZF0WW3PkJLmohEQUD0wFIIq618aSWeGbvo3vIU0OurB7N+JxBqf+O/yCzfDU0B/lYWL
kqn4NRmcDAsVS+EDmPw+msTDPPbV2cOsnFqmhCv8ens2YEse1aWtU0VeIZHsdN3/xbC6q1ds+1Gk
Sn5z91B9oNADdGF+/ABITR9xMuEcj2BV2x8MulHszNqIVsprOcgjiQm2t68rsOvPv0+j+yhJX3kC
CVT0UsADMv7lu2GoRTP7s2T3YXPW1B3oasE49PWCaqaQpyZh2EUzFQLOwYDIttJ4kven7YODygwq
qIyRMAm2ZK+Reo0sJvd/ubsaRgZJ0mzc1dOK15btejc7n9oXAMiLzuA1cmZfHrFijkGYSGTC39y2
+ptihQ/LlNNcsMJhW0ZgjgpV9/F8+w09JFamwvB8XsYQ1UB6GoLAA6qbATLouhmZCha59sU7rdWm
bYBpIppxGQRSXjIhDnCRQvQ4lqlHTdRDCrZLaNBQMRRRYkvQg1weq/1VUe01YfVaiGiPy4BUSTQe
ur2vxB+PsHYKfxA2nZwqit7vR4pmOuikpXMyhk/dliVMLTX+xEtNlSIVjun1Z7sJjMvd9wHm0qor
pMi+QFITL5g1Qp76v/TfNXHS+tcmyA1qd8rPgVv12fU9KAiXBFJQLxJWNkv0gUV5YM5bn9QgTA4O
yTRpo8wxloe73ODa2udQ9B8J8zvmYMnriXB50/RPX2p/8hZOmO59kUPolar4ui6QXZHfy/BceHe4
cNoJwNrVKry0RtHNxhjS04D2z1CnYUp+u+SJN2P8HNXgbjz0A+qpQg1nQ3TwNR4fzc4Xw2OW3M2t
OdRxR9cRXkplqemw6BRWna72KnrA5svzhFe9aq4OBhJ4154ZnLKB8EqTzJS5T6G+/HO7uCEjR1ZE
IyU6PLI1fLiQmtej/PmzXgWXjK7DukSP3Ao0JLutxypOh2yTiBzsbfCD0+GYT8UiAxZlIjhTcdVD
sRoezhvT6/+xEEIo/4Z5wdtiCy9/zOFdiJG1kY1/W/P7M5Zuz4NQFkmUasmQVitFfBg22mJabZKN
EJLiZbkQACPS5wqV/6HJkZidl0P2VqxjwY8YcuXFkZ8zbJP7s/O4EF9Gty8jp36I4MvU/UWGK/Al
PfPlWNp4670AAKBaQP47Kg6PdggjVuleUDSDErV4W58ZdR7+2ZSXRNknsMndluLBiQT0LcJ7Nb02
VjCBZimpBKgauMob6p+p41ghyAegrZ42q9ewLG8Xz/IpVksyGuwJbullmNuMETmr5XyGlzDYlf6O
yt0s/P2s/VrsxLAjfobQTL14/aUTW6V6ZSmYbD9xBwLZJv2SlAkJIb5bj3Lht+x0G5ZNpIbbsWVx
OXAHaR0vD2VYSS5vCix9RcTjkgjkDVuvx+Vvd8QEdC7vQ4TbilU30xAkHhthSQ3Jsp1DuptPpjOw
FS+fBYl8caIV9PKMNteBWTsrOxMFBmx6pOOvU1TpUrJyL6Lm8zkiOnJ8vVIcPUlTFeH4gLiKvElP
A28sOy+cf1Xamj004i5X0Yxe7QopGATMpbFk6vlMUIP8lA5qdAO0z03x8SD0VM//y1gaTEGNsbu5
QicyHNhu34P5zx6w4Cp2/zE9klf2+fPcQOdAiAKeG+DEgVvwLNRXRlEvqFWH/l8+AHPKi+6utq8m
VVTcfIIpdTStdgo93cSesWRUtADJxO+bIMg0x0PjcZ5DKHkhGc4J/18p1m3GeSVMNPrDR5rj5TOf
9cBNo8qOdUqZBnT/vL4yIKOtagdYnMmBV1BLrVvBk75TMI1T2jvFQJqWaC0VkQBa/YgRqHgA/xRj
FLh5XtVZd5XFZ5BalwNAvyX81eKL+fCJiDwpeuaOz2M3ayaF0F5Vl/Jp3Iv7IP+sio2/v/0rRHSh
MQM9Ko5tbBbOaCl0MXfgirYp9fVedVkUiZHVukpDrCF+nNLq+5QwVfLBfmKenfN3N9vvtBPeOBLb
6NTqHpRtV8LBZ0ZrqF7s+c1HaFjr1t3945QffwVq/LZNVJGtrUu/U94rb3WE39v9JGRwwBDXBs5M
iyWiBEUzMkjPpcFGQizjF1zbxSU6nMGjZ6OJFN7pwzs6dbXns7bq+Y8sASFAWcTIgHAKibtkh2wu
udAObYWWpNorsHTNaPFjJkpN2H9HGanOnYnhPvFQVfocGYylS12oNQAZy+bFkmYnwcWEh3KOwVpo
rDwlQjuhnsukjk1crizQFYu0Y5rTgHkYkrVVZu/jnC6MkLbsEYWiKsEVbmOQe8LlPJ28jnnnlnM0
sn/516htHON8uTyTTigAjjdCpjy5e1zd6GI95gD7wD8V60pSNQj4A70qJfdMuTNV+6LpKpaZxPja
KHX0Eso1Bpn3na6bvPny0T8SvS32L/LdBsqm0v/6O6NTYH+RtAfVGZLmAGJE8VzFKT4KJPmrkw+C
c9GI7teoE3WwVVMhBDhEPmCffPn73zyaOgobVBVBpt9W3ZvkUyH1Luly8+Z07iXy70dkTSyW6vK/
YVg5MXxfDKpfUxuYa1NS2UEXVlouRwFr1nNDaeUWU8XrIn74OY0KO7fZK5Bd2Za5N9vhBz9NCY0E
wmId6ftYz2k1qzLIucn7pn0iz3W0arqDzEPuO2RIiqFP/2MvuA/PPL+qZC/ZsFvnzqyzP+EWkSXn
zNc/5n4uWcnnBPAk5m83z+V9JDc4FhjwZwoc3rPICNxRcbQMQZG0jUMpyPE2M4wzeObQvCMTVUEU
ZNJw4uSFqzsIbpdyhNKSihFB1k53UZ9RwkEFQhpcwJETbbocst3x5SvSRk7kxmz55GJNydOFmt8j
byb0VU02RMEATUXB7Zs9eIsgC1dtEpcd7UjMpRwz4wE7MI9AM+lJ12IiqqnkzC1kQJfNGVXT1Azm
4zeZFe9GAdcv9yaCx9zP0vUql6nGAur5ykLgYEQeN/Uaj+Iekdd49nQKqlazgu/qfTKUnDCfjMcM
HXDykaCRWDdFcau4Fq2vhCV4eU5tgDWzNJKicFX1ewcTNpBaJjgGpr70F8ghMcjWSz6bJv1AS1iU
HN7HEMmVF0yvGTMwvwtBDHL4gd6Qn9+zD/5bDV40kE/RzADJNE6e4buuuEJmRtuX52wNUAofcB59
2SBikFC4V3wVBt4idZnTGEiwadiW+FFtzcD8VvABbG2SRRW8KLjO/0XGQzDt1GycsPQra1oGThWy
EktXHluxInMGgGgBsKrsvzU/MNHg8DHpMTy/ApphjKG9c9UslONgv2NxiWrWaNywMM1mWEnRnF20
oHinVY5jefP/qUaOKO6wtotySO1ARv3AxqgSziXN+8YmpFdxSXVENf7wLKjD0l5bJCiEfxZ+vvOq
0ahZj9e9voCinImuO3oume3F61mCkxJF5pdBFne6L/R3AslDW6JVmXlH7gz5Hbj2gi9eSnIhyobE
pN4SlsdEZyFhC54Yu+GWpB2tpWfoLGc2oKT2CWEt7qRp9gV52EI8tEPgL+aoGpzGABm9DwYaBQrx
K3xywWXMWGwYCLZaUUtq4//Z6PvfEepEkRIiktPKDWhCCJUsIpTf6zQkHkyz0VbDV6nw6f2SGrZw
mmZj+YyGv9rUoi8GEy8+P3p38sD5SnxMY7i+R1dGi4SMyFJCfDnAIUwrn/iHY94QXpbPRicRzIN1
Q4xbC3tsX/OitUu/cAPk8ZKfgmq1BK+FPwajdDDqrKC+TfdrV9mBrGE3bgaoCeF9loSoKHCS92Jh
2NT2DvGhW2wPdYpoWZwiLZEbuOFExJPeHy3W4CcEYHWPJGN996CQS6sJErjj91zmIZR6fj+i9Wlk
Vtzw0/96d9edn4TBqLWoU9eyjeYoCH23y6YS0tj0INux5q3jH81eaHgqpXwzxIwzhWbtDkB5uh1s
E8AUqAWR/gLXmj+4bIB+7Al59VTqyI+k3q9xBG5MqT7VD3ait77n862fGTIn1V0h3HnWdOe/ARW2
xMll+lMZcxQbYPtg105sa/uYXN72Hc0H8K7iJGy4e5hDkd62YxqOn8l3Sg/q8cEklM+ULjWOBlxB
S+th6j5frPa2mNV312UJVk5XK/yAftQsf8CoK7KbBQM3Ise2Pfg/WnJa66QBZwS36AaKyRsh5jTJ
4A0rE2oeE+akUDq+H5EhOYcOzU+jADq69bhoIUVRx/Gy6dBao34ipWBkyoLQt1rbTv9QGVFsZTyv
YID+BIBNaeOPI3RX1dMqRIpzIJE8q+P34lkwZ8rjdca5+FrwViPGzHzEo6skBfqkRcvXNmvRYfM5
SXN/qN045pK1ltSZuQtAaaz5uKYXWd+RNNn6PLoX3Jqs+XWmdbHxej8HUKVsM7D5xeab/HX5IdEq
UF/PzN1z+fwUxCyCQ4E0oUBV+8h30gA/oMzosHDATdkvXj9T/bAcVOJ1twHnopTC2MqpjY8XjYCq
USiBMC8Mj87TbnRhLCfMLBJ0YE99jGq6uzRhBqxQNpGhz15jK/y78j9iiULxzPWquBiz1VIouDFm
bM3MwBF6ysbdzLgXOdN65Gsp60USxbciVyvbnS5/65PgwyO8velqimDbkVhRAvSgdFJGnKqjetFe
712G0QCWdkLgwKYJRYT+JIYjA1h7nFs9H6YwlpRiI/Tt5HwiMqndrmVuWKhMHKuKALh62xzLOWBP
RkuzK8JL/4Xrg5eAZZskH16zArhOVrRTInOWrWkIUvazqaDVzwSU2X1eIU27cTZIzqt1RlaYpXT8
VVb8YAXoFdT09RUl3xyHNDzm6ZCcZLcH3SzAjZzPL2gfNZmmr69foamvQRGr5roR2mYF0YBPNip7
maevkFSOXpKzgJvlVgQ2Ro5br5Vf2oM94MeztAbQImMnNmMEWEIabovrOXkt1vhRxKNPlymnwG1p
KXF4Ym5v+1Qkgz4qdixYnebamiAvd3KAKfjJ6JQvAE9lrpr6tcTTZ6GRBC42imUIxj/fBh/2C6WQ
c9JVi+qRPyW4ABwCstVI3F5LbXsym/YW3B2BjbHPTQ2w8S91l6gLOGpM9Z0j6kmZCZHdJpsuaBCa
RmaksAbOvOdmGaEtWZMhwjvUmC7GVTWAGZC6xUXNlxodOMGyscdyCUnZJwtejqytb1WNxSMYIeiJ
+BpxNyDe6yOPbiNOr9IxGpNHevMaULp3s3PvMhlOOGijIDNqLMB+mM5+sxbHrJpPRoLORJXkujL4
YyPT8UrgeWiCrtiiPh0JYtqOIQfSaxLad23HJFZxddqv/gQO0JI6YhruF4uhXNvKC9/1FhUnGKTV
wrKdoiRKM+TwpkABe/V9zrtz+RNjJrwLWo7Lpzg9r4Mt+XbuQ6/G2wW1Ajb/s2/F5+UrqWsi0+fH
XEVQJHzkxA0/iKDNdElWvSRAkCM6pBs711msgZAyl2zrCMblvHuuy9xFQmudJtr5xJvkE9XOTvif
wKmESQgvqcUNLHiJuebFYB70JCL2tqrjXzXhE9B7nH3HOVbCU1jWsf4qLKbHxA5ZtXHEvStyLxIk
HnHeWuhYq9V6+qMzdOZgrS2i5wGlKsub+2Y+x16Fcq0Mt2gXNRQgbkQFh/IcypewS/MJldt5gXuY
qbotLdLkLj95+Ygmivap3rMMxixSSGIKxZuvPrr8dcIGtFJeYAEmL1E1kwccYJ0lnFPP8Szs5Z7j
bFX8O9UahSU1j6uS/ckhrUvkk1H2Qw/w2XtT2Zl+gFe/v3b6Mn8iCDyGRUbi4OaqWus00oQqskLT
STL3YwGhPwLehfGVbvQlu1SVrly8CvXa1HDR9Htnb0pM++6D9jfCxWkfpYulS2jus+3/uB089kJt
SojXHi1/vc3rB4d+jz+UTH5P5YiJWk6giQ0ZqK+UGG8VePHl/FcS02997LdL9qe90JcSCeCdnoHt
MYT6Q0yAKJBxkcVHhZ0wooEGd+gumyvRfFVfdl9yMCim7+kOX049EOl7+7gF4tlOgW2mX+Lf8LQj
rYTPwgXwk9brH5sjoCgN9MK0vnFl14kA8puSe0/J6cherSlTo9sxonU4tCNQkIsOzrCeY3KppF+A
qGcpe3AzyfAIqntiWLjIoGH2ZJlJwW/ykUiX+9p4JJP3/BwPGXycxB6IQ392abD118O/Phb7+DBo
zqsKFhOpi1nU2W1rG3WdryF2pQ8mtoM5FYHuUBhmGB3l0V9cgv16s2K271Hcp/1ihIGaH0t+KGdP
lzxuGm7nVB9bu9PVMr87VamEZoS6K0BFb2X34h/1iDZPfUHhKiXSIms8ZnSw9OAGTKBYR4OgRJY9
isn45hEgNA3AtdtFCnhIgkQYEItNdMrdCYXSWLoda6GbrI2Floo3CpTdRcz30Iue/lFDNJAZrm0M
vTT7kW8jIv/mOU9Tb2XqcoMUX7wrxjV91Rk89LcQ0QEJl5wOlrl7uWoE3S/5IpBgZ4VNG41ZV1rm
Mm+l1ik6ZQh5VqUmpZlvJoUyWv3S0ivHvc/qpIRhKrx7Ungqpz2SwIND6Uy2c2NhPfSk2gPvDrHZ
mt3EQ56XUUOsP/pmHSbqsuWkA2zXLZhHslvhZfqmCswLRDkGozwh/sMLjG+xZIN2Tib61RvNiCMD
+rLw1VTy3fIKS+zJ5n9DE6Kmc+0P15YDWrwGyVZw92j488G+Rl9Jl2hr/C6D7Tv3+ioFAEkcHETJ
ctvZV42r5JnJyNRQ4odTSyyYSlD17trQMTHrYDGh4OV11muvHOAvLJY2VHZGOM4+je4DC5hEfNME
wPySmsp4oMKOjZ+6EYR/FRH8cpJwM4D9RFDSBwyqdwvkft/TWEqrSFDAcApHYbKcWjoyVhfNRIZo
ko/+RqNjOxz6kADcErBpCiDxCvHd9fhXsP/+/7YzLenG8LPiS1Cdsw5JViz/8KQxoaH2CfqcK0n1
XvfZVLRFvtVYhDLRsLxy6x9or+o3IXKVDxqFYiWhYPbnwacXeLqWnXpm+EYWR5ySNPKnyZ/+xkxU
PS6Lb5aLWEVXAg5q5nqVMF3MiKqmLifQm+sOvSiVWBaT027CYWeMEpqI3C5jwFyLy3PHbst62YKn
UsEWxjHNdpRmlLwb0a0ASzCfW34ORwy4MdRY0YNTqwmG4/NDCH7SWPaGa2Nl/FoJ16wCB9vE7NwV
EWcVI2MD//HptQks+PjwGJWaXPF0ODjwOM6NdO0fnA2vhWEqymU9lHJujGKjbyD6z4mSvTmOdEqT
CzM3CZ5eMXgvMGbMkNLE55vIZRS+OT3t2DEB/RCFNaIy+BdjQDxEjXmq0/ZDgkPbGDPp3MDI+Adc
bMMHdpqy2qpHlgehM1HdTnktP2qWrjKcTxlW7Lp+joIQMzT9oRR8fvo16psSGs4U7dZ5Y8WA18HA
Rj5GXfDt4V6TlHdFBcoPfsCDdAHpIHamGRMpvQcmJzns0SfwNuv26ZmUrjQETkM78JHuCuOzwO6w
afTTpjsk1eIGHL6I0rfqnf5JRnlRZD7U9+r4k1EckiySPxfE9upiNYp3ujsBku6wFpgM9yJewI+O
tNxXJ1ruCsorclTWuRf9nOXFygVTx9T+qC/8eMpygDgMiYrKc2wbguiTw8zyAeGZzuAThInqYf/0
bXmhUEgIuhjDZqhzJmzUeUSK3h3MbgbRRIydvw/HBqZP3+24XTraa6xB0iiFAxR2YX1lJmYH/qVm
RVKO5DUfDZg/z17jR6W10kzRmxQbHEYmaE/LSFOTvgHIN1ig8wKqE6TD0noQuxr7RKFh9gH86Rc4
EOJRL7Vw7PquZPSP2BsvrieW4vFaVqi/shF5MGZJy4QSODmj2wyJX/1ta0rCMDxPMDIl/J/bXO9f
RqcBENBjMHLYan6fut2NiBvz71tP7wglBY8cdnjqYnVlNWC5o3+EvAdxFa8apCy0Y2tAVzKFw4Ba
LqceZlEqd74l6ZjFMMG7aHnWtzm9USW/4Um4HVvMUeT/7G839quZHIBdd+VuPBPRvHUh+Ostlt9h
brhYh0y60Uz2dZrzG7QMUKAQQHwuCVUhWKGq5mIsuy6nZzqjRKLx2z8Zaczw5pcmwel8KNapQ0AJ
ZSxIRb4ZCQew+Bd0eMyawKWyMvipC4Q16QkIdwKoYN3lrQrIav4LS4Zl8ng4TFKk9RkyOHvtt6rQ
gBMSwXmAA3udYL2+yNgLt0/1SSmnPhIw2lzV61Ehxt3s+X/OcgDXOSMTa1IXjDgbEiK9C9dI/drt
RGr3EVb7PwhfqOVWF4/yOlZKOmbAUPLIcad5H+ODVx3mcFFUtAGLV01O2DGN5rH55gpo1zoNkTp6
i4HNgPTtpJgKBvA3BdjAV6qLOXJVkGPbkbhEuTl2R5FPu+3D7O+uferrxxkMaBkhTRbgIAze//hr
stPcVZYW6g3tzPAcAUx/1KJKH1WKrUuKlfSi2MV4roOaUmeMVA6pTVY90SOHeR2dfy/KMiwk4A0X
jNYzeZcqAmNMr/WkX8VOeXdUtY1Hc3hUxgblVTYQ1VcCLyAYrnSP4YK0f2ODh4Ckt3AyZ+kTYCNg
UpyWZFhOX6G6e6X/ex93rhJm8bpzc8O+/z0ZOnUn5vtZJT69oEAAgTJnDVp8zgyxr1MALVsXClP/
/x8UeMAg/Gc2z/7hhc6JMfADWfalnlETrlKpamE9c07UXJxgVHrEqWoXf6zFLP2YKzizbt3SEsnM
ojK43SevcJDADK+FOc4pZYThALP5ROMp9jzkxLOvrVXut0q4OEvzN9sTb8yUXGh5lOlY3maRJAeD
FuEEwDMs9UeHFRrRy6pRhUiw5Y2zu6Ds7O52YDB7c1mWwEDEgq9pfOsrszmiZ9ul+CabN+tfy35D
+NliTR10vbDFDJdQed7pPQAcBh3HH5uC5Hu2nbBtgZirwuX3NdzvXepWpFJ5fScZxRkoXItJXG3D
8+gHu0pH+1+b7o/3IJTPYxPseZINrejy/9BSsjXspiQ05c4tjOS9q2pA6xPeW21KUYW9kfSHsgro
v3DVNBAV/UWrhXKr5s6ylZJEpZrr0mbnu12lSDGdPw6Fl27YMuLDr0abLLzhrTHo4Aa/LCKOokD9
ao8x5CSQyC8pz1KTnZLMk7ZKzHNbRpn75UkDamsjWRRUDEDnIgNURTg09lnMJQ/BkWabfIZHfdHP
6I8GiznpP+gNTt8iRZCk7MS1hfvtvm6WNham3G9OfAs2ZhGJFWsTuunsisZWSt6/joY0Ol0c4dvI
09Ozy9zZiLPxn1zKiZdFe363f8279meHQFP7rSQxskNuqh7pjYeZHcrOTJwPb5DGLkOWzGFQC9XN
DHBOaLQgt8R609FW27WrZe8yR3ToilkbObAlaUP65aRhxyXMGwr0e/v7Qv6LeeFR9UZhWYtbfXb7
YIt7NjgoFhYKTMQ5z1T5TzbLttVXZbjDVhzEiPT7KH8hJ2STVnbk3cRMpTlQ7FGgvoxY1BnJNc9d
aV7j2eAzqKHu71Z+TEVlg9Xhkeycmo6X/v3MMkLT/xUzfpFtyyXLsGriJV6jL9yHHK6Fp2F6bGJR
TQuxjBGeuGssEQ+3e/AqsvETJNO/ZMKWsr9IWGBXC4yySdabcP1p6Yrm7YBCX4VOLRD0pn5rQlhj
EZaP4xvdLq1nmhvO1mwanRV7aRn6GLx6MguC/tK5EY0l5s5Zv/0kO+i0LEbnxN3JrBi4CtEbaw8B
n68hdn24wzvvzLaofAuSYu93TmowxWGSu2CxGuHX4ZPYb7HE1fCSiDLM7wbpLGgFilOOzHC3f9/k
ybFdwJ6rXUaQ5azEs7bUNQH1qHr+b67YFdDHpCMsRN2yQRnLuWPJYpCAP8jW5pEWkwMJPZjxmWGa
RUYYEK+O8Jr8gigNNuhm+RtEI2J3t6LjQvHFJz74CmlebhVrHt9w6M4cB0knv9kwve4b/uJ+tDao
Xgh2QKu0s+sS68I823IPJ1OyRoNDQkTgrpFvUEJ//EtPmDfdKjpJU4qZ8w8ijwvWSPi+CNYM7NTt
/GYGegawKqK3RWNTUuIMnNAcZ6xUcJWqvujPbaCg60bNOEcKat/EieyHRMZbumCrZSHrLWDwA3dj
vyNtXadlVWZ4N9JIUd/2E7Hzpn4BDP2RMug4ZB1rWjuQ7yUIwmXrJO7R/+SzupIjtvug3Ke6Prpl
Yooue4Bo0W+yGvmQYMBmjPwbswpzMVlkv5GltxJG7JgOLiXJJt2Oi8vTOXuAYbuAsc0KFOtf6Hqy
xgRPP9OtOb8VTQPfukur0EKrdeE8gHDxTWK+n/j06KRvNJZ5RwJwMjJL+4cO/wkPEG+xM7x+YDc5
a+1awV0/xF0FRvI+dOIoGR0CNir6QEeMCPQEHJvA1pXsE73jWjBvdvQ4H1u4AX7osSVy+lU4r7Os
JYWBVIUN04Wsr4tHafKW0QQaTf8zveri5hv/WaIwTY6rqRakBprMH6Via4Mq+m7csrOC70Fe1XiK
vLU3i0N2pa0RyR4/n+bncdWm6FROHVXBsIaR7BYG8dmLXi1gUwmWJxKUWLNHB3UkdPo3UhSfouOO
3/+8nQXRTbXXq/e1oXw+ReTGoryhT83voPCUQNOSBBRVJ0gOCnhNVYDl+TgEYJDcAg+3yuoCs6O3
DGMKVVxgh5DfBWdTXmoYcHZFM2yHS2Sl3jQCa7BamM8bNFmAJjJOuJLQK19PPcO1jTdBSX66r2vu
Bd4pmONUl2hfCrp+I0Up7goKFLLtEOP0bpXVKgmySrKRCEZRxAuh/hybM/xlf5Ihxa5FGqkAPVmY
LSSbZGSHPwbYObfGJALTA+Bh/IluGCRrSymg/Lmv/tLPRWVrKyAPG/TCkllIK+qLLRBseA9Ve5ma
+WZDNuJUuuRnKLQBAaQxpLoUxvViqlHT1u2bSetukqlQLllMg+If8VjaCU6irT0az3fKhQ4M4ZfA
mMilRKlfeTnzaSlHtRV5hOAajvg2VTVKT0+hhCIls2ieqOjhLWx2mPe0UYlNGnVm3kbmnFo8uw+C
7hHOdpIsdq4pVQbfd360DJvA/ozV2NAtgNvjn4o8MHXUQlie68r1nVLiBit6PX+VABNM1dlt8ME+
YOqzKq8c3YUUPSZqW0ny+G2YBRSWrYQmgMnCHGjRJ0sMef1dKcldMBrvpSKKYMC/c8RMKjZvSYdl
r1A5YM+LOLRjvJ66NSVg/6bZl6YAkEh9OQ3Y8pJtKzy2Oc2Bt9NNNOliG9zuPHB04vxrLHeyIS63
s2FnI/HeEA/7MDPI4ZzxNNbRVayMSvniUdcKdBAcGKOSB0kSPW5QFXJ/3BcBox+iRMQND6bxGUAM
p6r0bxS8Klu0RTSuiyDt5qjDstlSCg7JnKczIK5BlCo8RYgW3uMD5krgUYUAUDt83xLi352h+JQv
Gu4NmZ8DQKgrv6UoauGBXLYy7MoGvCCi1GAyXp5SMazCEy7c7GS6tuhlgXxTBBThzInM3c/w4WLm
FtsnGW7e0qxxnzFAiL/M0ybfVj3hAzcxWq4R/WNrd2MtNcylF1oLrgUwA49PeOwZIQA8wmBq4Wrz
K2ocpsu6/MwanGHGAcT+MW37MHN5hrdDcwaKCzoDdb6jTfZMLjmMLxVN/B7Z+C1XCaXoS5U4f1FA
hubuEom/2Pni0yyRqWlPolTcfo9DJyv8llGI1oLMXKsuRwdf43JyufurNjwfmx8carYXb6rfmFuQ
gpsQezJdJZ48MGI/XjX8WmgpnIwi4zpTM9+hUXD+U5AboLqQ4XjokLTakzTuqZjWjxvVEsq5GLxt
AsjIJ6jTab2HMfLgaGGh5kEZBmyJDDTMTmxC0OqD0/Z/xdnKF95T6iEaXz1cTXSh/vIR5t415MTY
KXqpmTZ4Hf/1qKg8NP16wLjJZItKrcYns0Z7mwPHD/mfyLW5UrlESdCt+5L+AFJbSFx8QLYhBh5E
1VG2SKsjG01vn123DeR3/WbRBHC7XTPXug6Oh9S3z/J8Gt9Z6nkBToM5VKFRrtxajoCnlgrs/lCQ
JrXti2YyApq7n2yCJhvR7JTdAQVR10jBGBE9X028MXKLZxcTiiwWxUMC46ESg8MireFatmLVUJds
IVIsg6tgAXCpgiBM2C24Dh1qJU0Y6Nq2VHpYJdLs/CO21Fvratm1mYBJxsZjzVDq1eTMIAfA6eJN
3wcOx2PSDVV/h2VdfCY+mT9iaIYFREtXo8uWvVUjM17fwVKgf7X0njmBlTWcgZpm+rLbZekOtC8C
3HXkA1qToQvzq5oKBDTjFKiZIUtzOl41/MBr64e7N1qaM9OkzjsGAhDrZboZbk7KR3QyoDcjYfkI
nfxOPvycr4p2owMbI4lqmc97FLB9PXXT7eirCVXncEYvvmAUFpujg3EwACP3g4omA0lZ+WrWxU5N
ZUG+U3VzHxQSYlYZyBmHks7twi9YtiL1vNQZvLLo4xkj6uWLqB2OMnwNfIFatkZjs/8bcym1xt66
SC6np8tl6naG73xuNg7oYP4R5X8cqryYOEYMeCJqWh0pJUL2QpTfAq0edEQGdvLLw6eavotoqDe8
RyNgaBhmgiXywL6LYabGcOxAhS4rTkhsImIqRt3mKUe65AUQfWVAksTfFjshsYWzyr4rQSMGE3R0
FWB5JxqANQ3sr2aTTbJTRX2hHWax8k9lI2uh/PDQpUyI52iKaatnc2x3k3b6PgQlned6xoIxxvab
4K1hXLGZldC1Y6knJ/epKC7rJVBYWq8izgvUayOlCgJ+iv3B0apG9DDhmSLsBSaxJNXYnK4kNGeH
wiYqf7050dVFrnnebmbDm4K57jvgmmxTVGxBZIM0IUb2FaIaKlXxWcKumX7v7/wKI8KxaMZNbTD6
zQGHcXZYkhcgFnPhCV06lBO10QZ9YSjtBBclLvw/hscSTwCy5eKksEVTaAe/HMPL309NQRWAzuNe
X9b2liOgyL1TEw/riGs936dFDok4l9VLhMq6tJqrEqVrty4Ka90lshXbLhI2+dc4hiKKB7/IacV+
LcDwG0larBzsHQir3eypFer+4bErA+sCkn7cYPzMUrDmxAtHjG3oXr6elUHkvmTG7hHBd+gObad6
OlBp1uVOtUSzpXl3MP7MWp9FiGcybWrVUU9QULQfoLxcgTZtyQkxyjSiA6po8czqAOpKL/1LbJDr
/C6pl8NCDMLb5AxLbA0/GnNDmw7V6dU4J7XbHmx05ppeFjEvLc9nSrMcpcLJRQ5UktUqDryKeftE
W0Q33h3CXJMOVrjh3NbPXj519nrrLnCn5x49OcRcpITe3loPOgmG/opE19z70c9Ug96Mqoe4iOBr
IFQMP7juTMm1r3Jj9fEfhHNrdtfeaJcZb8JjzPoIh1vHTRM5S9wPLGnQ4n/U0gJX0nC80N9hrCAC
fRceJmdtsw/aH9hFqJpy2Ry63uXEheliq5YJ7UA/KqjtvzrWwSCALGXEzSLxrq/lCHB5uVs1AT+d
j7+LdUDDwcvfulqlN+x5DnGgxoV9alcsqVhD2Cj1ja4Qq2U89GHSVJd/UZMZCK4kuHNpisySGjFn
nT45I0JPJSUT+CUz5jHTUH0/NGmwTRXOynYz/GGWLZJCQZUlPdn/FaElxXsdhb3FQgk0j2Ov9xxm
rA2Axgm2ixRf50utuvuMAj2KWYTylRPTLho1payoBaVWhgsakmjil1rqASAB6kBqF7cy+9HfPktO
xaYZB3BEEpZcqV38EuuZCt2+3e9Uh9TI8i+R0+uLnioE6deIFNktGpiOcOQjGcCcSSOWIwQDul/0
0C/RGFEMJLydocpAzoQeAZJ+4u94n6wI+j6i8XFuX075TWla5g1uDP7hZ2SlrClSbTV1uZstc74Y
5k35R3u1lxmdwJt7JUFVOB+X4ga+LOMlwQuiErotixjypTtmqNst9NWB6Bh7nTuvNK8bEEEoG9Jo
uJeA+00xyp1knRvoVvtKtaKzMAyt3ryw0BEizasGyYgQipqJsfWQWuLDmDimgbV/NFhQG3CgVPSB
RjfkbVwcO52UUL/vy/ThHHyRpl/OWzGJ9k8dhaRsvAxWdRFMm2l5OTLAt/XZhu+PqNIrpMjh9M9U
nytEy38dWBx2BEa7F5RXFObhw5/rCRXNcDuugJkdOBZvHByOW7MCq0u5b7ZRrpj2Htx6Xup/r2V2
Gly5DuDLDzBwkBcFcOhRVzrdEjGIM9V41AhZ403JYG5UFOC9jM7yHTbWfa99kCBSnJY11m8xUHbh
+t9+FylMY9ufvRI12Xy9tmt04x+CWjgds4t9wZ0IguHzXo2UL9YSHuyxy1RbrO0sRdKnNXFmA2ww
OCV9U1ljid9modxwu0n6IvKBcgjyJMP55L9o3yAeIA0fMRgQ8OYESLxbIrx+hmJjiX6wGLRB4i/K
wSOUmcVh7Yv1wJCYVgp/hF2PGcp4j0qTInOryrSaldTydLL4+bToHZdPraqeAX+Q+tQ/sGYAnix0
wq8a0JbmMqtbTxQZCyi+t2bphXCArQZ81KN3qMh8urcwxy8H/yBzCghWK6EF3XZXT/aB+KHmo6/x
XAMujXxKhHQJ9OJSpIkvvFPXysiVqtSObCCHHcKIF7Os85K/J5MP2rR0/+aP8Pk+LMQ+hKrNpMAt
PeWUl+HNcYcR6rbCqJMMa0foDFQPktsDHPhEPT5SUSl25Ve9dOLoTJIi3fYj8SyYu7mkVQ6ZFWlz
eroPJEwlQGQ46TypB4RY/n/6HrHfJj2H+oDTC7hOcIvxoetnKbZprqvgbfahG128gN6NFXVbgTT+
12SvYmXKCV4vKkZwC06rE53+HrISTsHUxs/YOeOlr/mvBfmiEahvqjHay30BVhIjT1aHjOshY/Rd
5WQ/ON4HzBH1FmgWX6QkV+sAmWR7K3P7lt/oDNSQDlnV/KlByZi0gAq+P+ppkzioyAtuL4ipPrnu
xAmpSylSpB+ElwwSy3Pjn+swYvngzX/+pD31L77BcsSJqhK4311M4daOAlRdVnzSIKExfUV9sMJm
OfXj9R17l/b7hkFGTLJiyPeRhs7iOdC7i5C5pqKySFd+s/IPnNJ8t9HoxvSrQd5YzM0IcUkJiHDc
m88tzcaqZxjH+grTwtXyzM8DK0Khovwc383A1LVsXNxItQ8vGNFatr8zE89D4fWRSMeZ3j66n9re
2AOPxcnHlfR3dOJBYM1lrWR1yYFu3eBYeB3gvijFSZDOi0xxylf3Ope0aqMeqpgTAWvwsUZjbGxE
fzXkyBPzGr5pVCGkWNRWUPq6x2YgPm3wky64h4oiLlI819ATmdpelYU6C8BAd1EyocraIueuyCC1
74toQ/GgkodgfKB83hWP+xHAtf0EjvQ8nyYrmH2uxT1Pl2y3hor/Los+QibqaUK7J35ITgrFv83J
6uvLCLl9hohOj6lA0T1GeGOoZrKULV/C0+UJ/WderWWw+ahmKwn7UmvLxJoYzVPhJu62MWLGfcZD
Bs4fJ1WtH/2Ov9V4Rm2Qku1hoyZBSUlCWFi+UXWb3jNIrnreAbmaAZoO277Xcfh93hl7nABiko5p
2VV/to2KK0simiCDUufm4dHS9bOlyXnc8gQqlpiDqQpOVaR4glc7CKiJt0Ir9rZJRMRnsUx3ZfFz
bvd5df4JIkJCn6KUOyaW6YwfO/gZCwArV/UlOEMu1BZFdgRuJBupdgpuX8TIJCZZXUPD8ccFBkSe
lJ/sODEclEd/BCyRNf1THqfFQCpSkH1Unz/0qFS2vO77Pk9jWfvYLl3Tscuepwm4MC94IiKKID4q
QW2jwkaYLdrTCZc0IkfZKYW8x1MWa0BaTUmM65NAk5Yo1sERmAMJ3H3JzEpWyvQChr4larnPMTUb
IvVqkChkh1LDwHwl+FUegSO+9pdZ98g/66A9LD03CKdB54G0WSMKZ1abnaSjwcRf3ClLsDfWbWf3
FDiKVn9L5Y+XxnDLtYvD5KFNj31XMf9AG+hzpNaRFfaZcsThoKdG0CM79Ee2nw/4S6xyB/JxSXnM
Tc9ufEzHGlEWbVg00o7jO67U/EVhnSfvC7a5O+t5v7dIzcuJuPgbQqQXeeTOsHaYR8b1tl5Gibfy
XKPrQwlc3akVc/bMlyEKoxPI/mLPSf6+Pmq/krmOzjTe0flbjEdi/0f0y1viJ9DsXdNz63fFa2r2
QAGf07CPey/7OBrn7VBT0jERlx6ojATDmyJuCRu0DOnfDFZALO14Izc5zV2U6zC/D3qnDilIMinC
PWsD55NvsOWcis2hldKaLbWN3UQnk2AZXWH/AOoI+MTvyqU0cUEBSiVuwYsoodRzbUnEa4KBQgS2
J/L5cKtYUJbbNd7pIpGvaPXIG8aLcn/ECKuHyWaSSNfFSVBHfyU4H3xKJakjuJcVj/TorKsxLRqV
z/XqmuokWUEoiGy+NtS8AXxsNURlCuUN95Knlz8Vo6wh7PRNHcfLc0Q9x6DtATx3csS+Ofo4Vnx5
itS1sI4cc3XuPUHNo5kb/DqRtKmfkS7JhlYxEGUMqiGwIaaiWCxWEAydCttO7hETWLJsJXBIbMVF
JAZVKqdm3x62htC9keLzSFmNWjLKtlUKFgHVyx9G3ZI2TiBIdr9zki4zPSb9v4sLQxWswBgw52Rs
Y8FkcVQ6hqFb4pakGCEicvqTHPOndqLlgfphmvltRU1Ax+prUN5pptHy8SecSYYd841SF8nQzPSO
gt3PV0ifrFf38Y3fxbDc32WMo++Ew76bX4lGEmOZXj+uLjm+DkAZWheo+550yoNlpfrqT97D+Jwg
bdR6GCQhZYRm8waMQFJKCmp6M6MEt5bXl9dtGsB+9syDcVd36jR97arJgK7SN6CDB6gxkZw6cbT3
qD31E73hdY+QJX0f11oKxnr1+iMitkdBk97mjkDczB9/EV5AwW9RfdjpUSbePwgH+v3YvNHo1eRd
Z1/+RQqehCBEMQrv88L9oMCeS+D5WsBCQObdTqhhIubElEodGmEWr2hJqMDm9dL6r6wwwU6ngfvj
GFSnyA4S32dItnUYfkwi4rO9H0TlWXmS/EOiDxfrE/3MWZ7CKKB8ATLhIs/ZgbBexdxFhqgxQuan
D4EJ00UP8Xd9jQYr+39buHIOXD6bRujWO39vfEPhC4zKNTOC/2yGTOCnSDokkoszZvL4MkoYRKOL
Kni02hBWlxZDfCOwHhqTXm/DctOfO6IHTKJ5i8QzbNEaHEoeDUQI4EJtPYueSQBUMHZcp5PdB3Jy
KlS4jbvowb3uMs/bUhoiYYR3vRol+Xy6QtjSFuiPIWbdsly2Gx4GdD13gNPq/EjlHhHzWlAnHJM5
xK9KyTU711q7ahS1KSbzkn0IcfUr84kXHpAI+isVnWh5XOr0394LvHxRRHIzvmdTLsgM8/7CUfGw
wv1ABiOSyYMY82C4eotNLZSuJmmAFOiu0FikSTYAqV/uSgnaSPJnTvfAjs9tUpWowe6MFrYCVA6c
zpS8hsv0AnpXibA7ZuGaZA5xVqaDznh2gYb/ExRtjS6KISRstP+GMuL4Qduk4A7Jbse9MZ0CQnjv
rv2Q8pl3RgtZcINuTd6Qn3w8ReBtotHM2X+017H5C0vcnHicz/sYfORjvLh2DgeqoPsC5VlewhXB
+1p0jkCq5Y1TgEHdCEVnzJhlhNhVUypGWJOguhPPHsfxu0e13aivfTumogwf1mmlcrufgiXy4HFG
rJN1B0j5smE2JVauv/NetcM3woO8POMeXLeKpbcgxu5t/igXdVarLJIK/ePOu4haQOKjIB/hQYDX
De1BfYvkiTfQX73yjPx6ZxRVbxBAqffqsXHA6nIO2p6etFLg9zqNWZDZQoG21AarFuxjhIfTvAv9
l2mBoLrCKD83e3Ej8leaTAznnEc8bIT3Dn1ZCwCuxDsfTvxkbhb3UZUx37si935OMTgxQFGZTeg+
DHkAQ2z5JNQIS1cq6hvmpUBNkViIvGIpCXfQLp9uhOFGGGTrV84cCPNuGfFiuqc87xHGSFN+d9In
tj2FBtvhN2jzBH5Pg1lwfj8MhRNi1kydWd7ZbPW7FgSUBdhXHUnHfAg5pRwimwMI5VKUnqbXATVf
zh+RyX3hHHSB2muq23Mq1T7GLzwfBAcOAQeNh7roebXr6+eVxej95FptZPSgaGJ4f5MSGLvLo/5K
iFKkCe3MnkvqhV/LJb39Ob+du/lLM7xwDi8KuJwgVUYq3c9qla6tltdTdjI8S908GqwQEYxBH5Lh
2gnCZMhJRMDI5D4sq2bIPoM090PH+/Se+1NSsBggf+PtxF7x0wilSDROA1sg4c9rVPEUp8segTO0
AmL9bn9qCadoc9ymeClbPcA0opjkFoPcHu/pKV23ssgRRo5fPeCknosX0zPxbvvItuJr8SYXObJX
3RPUYaBEsSjCm43tqWPLKZ+1SQ4Va3DgxzhHIHTlHj1vOHY1E8odQmdI+DOsGgMJkqJ3clXCtVga
uOQROrM0E2gpqqKeZL3EhDQ5CaInfLfstB1eBTBQHJ7unEJ4Apsy+TLZWmKicdwnb0FQFnsgiVe1
4BjiEf6osp6Tepows516t8dgVaxQtS6cGhIuDK3HNphEuNOBN2Up4LrvJtlJ1kzkmfnG1/YAjGOm
RqPjHtpfwiOyqqXhjFAsI/NPxwAa1KmYj7o/LEPK0KNqpDjIvnZoFWOSxOgsqHlHthkkHJvjvNfA
nMgQeskPL8/8N+Ha7k2BFpTAThhFFoH43paxoqwaGXyS6qFc3iDBK5mUr3sQNjFMH2v7O91kWn6z
Y3srSvp8h9wZoXwxsJxGPtuDmXln9OT8F2ZmN2gk6yEffDc0976kf8aj0FmOY5nGQ2CRVKFRfzDQ
7D7lyCPftEdh8djTsThypYxkPceH68IfjZGRvPRYU6sEZVu2pcNkCRxQxvq8kq7S1qBMpTjrBrAJ
2iG3494WZPA70hSSHoo2PqFVSvs0KpHqkt09gO3ndd3E8jm+jJrXulTAD7TfhbRT0G/8MqTyN9NG
3moIiDrdiJiOaEyJEWA0bVsuzw6G3PmU9+YTLRpdmauSsMjtrUUFcBqS8wM2AqGr3uMl7webgdX+
RXqeoApihipTQiSbx2GDpox52zaZhvUACZumOOqbwwEfStv/uIt9m8SbJKicji4rm63GoFA/HxdP
lgXdPrAx0L00Sg/B2BVAuST7nNt+wFTtt19DxLYLGq0bC/YIQjxceGZq6V9GSBhPkB+BekJU0OzA
4tGhsMzcpL2ScxP/4Me19QbqyV4rcC1Us80NQwtSYUQufXOljZXEel3u0ExwEmiaMb+MkuFyEQnm
3haN04mK8DvT35H2jP+NR2pSGW1Vntc738/WlJSTcSmK8mc2jWp76Cc8mVUGJJCm7PuLYJjsybdM
cT26WPqQODrEUaDH3Dou0UKjcyajbFUNrqJbQBmrrTBo4Oy/DlTCCpUlgSN1sN+V19tW2z41CthR
TgYdHHEhDVFqTiu+Bx4rJUsOnM+ooZSqWghzqkS4uH3PLLyEmAiHqbdZB0Z0Sqo+LrJ7Ug0o/jMh
OwtvZH/U/OcUX1VSJ7uIjRk38DYgpUBrtQgDJs8ygPmsdgE4N6zCIpisXFHbZjwgMAVLuvpgimTe
blgXd3GLmwqj8r5KPbc6XD12EqpifxQfMW+sEWqzpAjhUtcm4GhqzC7Y/IE9bii0rw8trRYLTXVE
1hcJutEo2zbrMfrKJmQu0FM985biXNrpXqVfgXeUNiXFV2NEf+zn6igx467yl42f/0ApVRZDvagt
OioYqAY1NihGy+85s8c0pJ362mykYdDNR3U/qGiqAHXhQFNsXiDR4ijlin0AKhLr6jktYpeXcWXp
5xDwLWgWQsOQqtQ++1sU2lzz7+CbPu0b1uzcqke/K/exkWRVZA1CdH6A6COjNxczE3psqSeQ2nNU
T4s2BFotSKrcuFmIqG14fPYlEOhEiCIRKn7ZdCRKNL3EAYROJa6QgR8MUYBETVxdH3A2hd449Ypp
Q29oKfWM5VW68JPG8WB7fUPAIdHby4AMKKn9EaJkDcNd5tgru1vLZ7k8E1/xQHGS0A7Mmh+y+OyI
mwYqC4xcDRtHlXuu0OtURmvxbV1Blk+iA+bVWWE4j8uVDcPo4fBevxOzd8UJfvugVGbrwaFmPN3r
fXXYnCi4x6KudxF3LsLgWLM2rxW7P94rMW0uTlp+uW/FRXGfL3fust80p3x9uG9ek4rsRYIJ89HY
ZZe6muRE8KMGaQiwVt0Jyta/Fp7u4lwKA5Z0+vJ/SzH/5pYf6bVPKpbUAd9GgkoCla7aaCMLeGnN
7L9Fx4yn7jzReyCDeXult62k5SnWYp+W7IEtDKn8K6jeW6FuNK6QFg77BOp/YgAzsiBzDpsPl13a
vY4yXNd3Uwv8MQpW/PeEUVGjxCQT2zwCVDyhUsNGnBmOkfGdN9gmSTYcogLY611if6/wd4/sIJKI
D+cu55dQG+jP47GT/LlDsXlT7Su0BypDBroAs27lH/2ngcVWZBpjeWgWoGO+/3Wkm95l3QuUt0FS
rjFMn6ckbqXg1DZReI6PdF71qmShzi/xF/iWvk8MPRaeRcJhQNUIBlIgaFnc2UrUjZpZfwImo6jY
/x9BJtj8FzclM44W2aOmLH7pcKW0elX5ASuev1Exm1l/e2pipep5jcaKOaZEWflYembP3y1kNHL5
gmDpO6KEx61lir/3JKqQLI4A2TS6dYKOxkMF4mn0AfPGsYmpI2weqrwsKd5bN4UaEel+vxKXL466
63oQ7ylnrTKFdZK6n+0m6ZnfwpSNd3yI0YjmO27ThV2seFhgSCSW+3PhwJQdlU1Z9lpqaBg4RrIK
Q5kWclAamm/fi9Ep+M9adtvqSnBFoHT79RjCh9gaSqArri4gYgqANOuCvRCStVudh36UaNPv0c99
bu6UHqNDLSvpqSsfKeFLOqGtDsmWpyiRHcfLA6DO26V94r46wgYQgqLcuUx0SGp+Pwe06apWi71H
VrNdUaR9L/ZDMKmE1z8X3Eoyf+HYqg43TcgNXrSBn9HeeIuZElpbJJoURKUeVy6i8/grpNgWwBGH
csXy9VWkJ+6xc7m/tAErYowwZ55Qi4QRV0LMJ/ivUhZkKd6yqhGAak7jxd0ic91YAe9ts3ZUOPhb
RHfTrNtzfNLPnAcKHpdGL+vKHHzTWjA36b6uS+4qX9jdLvX2J/GP6VMxu7YrBqq4Ox1oOzIRVPFB
RzI6J2zfxa5dB2qw80NwyELzJTUM8VckdFZNt8uUTClk3kMzFXzOtvQO7e5P8wdgdjQ5SWJS4AcK
6sI7YhaHez3dNYjoUkRb+B6LGHs4tgLF8yrZ1PhYwi7sCksygKS5EzYBZ8Ye/s2m7i88saaLG8sP
jndNaK5/+hajCmQvvATh+wkY3Gl48/AtdqM8KDwNqLEqBeTb5FG3AZouL5iJumHf90j14evoiLME
TdQV9cUgw4CfukzzMmgg/be0FvTYaIgMg5PuG+33IIlpweRS+Be96qZsXsMa5E/RBOGorgsoPxRU
WwOkU4DXTMS+Pe4UhNu5alYXFJ4a5PIgtkNTdVys5z3CZm2e6Qf64VUv+0cxQgE0NGa1bLhmxDvd
gS/GO3Kwe6nOuqxeFTfl+R5Vr6Uic++/L/DFExb4+8v08lqBzxfwZJAAyO79zV6MAt6gWHwmrKuI
Zn29Bv5hMzb+3Sq8JTbCPuHe0qF4DO+/Lh3QrdHNLzwAHLPmZpFJQMY7o9p6GxT97RoFn51Vj288
GHOHX4Y+lAvHtVlKrcJJgbKK5ydrjoVlIw5Lg8wy3cjsIRrcvakKcYMXJCDkELlQIbiaTXQT54Lg
dIxBQ9ZaVJ/9y0p7fqHL5HkweZ8kjnW3/yCYSia6c775Y4rSI2gk8LbsM2KRRZeKDqhukLs4VfEw
T3rhiSNhARlDkHKE3SVBOWuqV0X8t6ByP3sweyYggq/bZv+3jR8fZQCBfo/qsG+OcIThuLUbPLKv
VSUVrmODQIia+Lari94bhX2w8YiSncDpO+Q931qcfUnBBVOfkptmzyGFfyLJj1+MbNoWtFu+IYAc
6PiraXUbkTGuDcviSvTKcbEH/7IwbyYMbVw58gcWmtedx6XHLUJSD7/OAv+W1f/FItzcpIQgkfLV
xMfmgZibhqBMPTsG/h2LbYLISQ7jZX/gpo1FdPlTIZvMTNNKl6kA/xuOZPVVeGevR5vCMMze7VDb
frFoH8bJPzqgjplka5IthYJBiMIlxEYQ30hpT6bMbuT8TQqIf7wbQYZUJ64KlYvw8lXhbAC31tHp
Vox8460qIJ2LqScjukK759+kzxymUY+MMGmvKkdwdgoLg3DnCz0c62m5bo2qhfGr5VnheSz5Sae+
LM1uSSfV6gTUkmRAw4UucI9/hleGEqA1Gj+whZxsFbH6WngrHYvpPH5ri66ZcnVNYFiRCAmGViFY
UnIhIi2TQnKlbMv6X+VNO7K1/mjte3iRtvHTaybNDuQEZz4TslzIuvNGLC7iOBpY328F3nIAhadX
AgcQbDXaIFnojKQPXVN6MEfjjJHYfholZpKVaA2mvVaBSps/B6O/Z59cpI56MZ8A85KkOW0ugrEM
5GPNRHa5eP5cgtv5kCEZPqBtvbnGFQXgW4YBgX5KbxvxHf1hfpH26TWQlSARcY09M6TT7Pj1H25O
ZRYvudEbrLq22XSph3Vkkp9Hb+D4jWHK00CkWTSDCaN0nZoaOBcD7yz2xqeX2nneACx2L94uEp+P
OWqDVcEXxzBGU1JpBdC7x//h7GFQgknk3llbu40vqHHST8wRYn7AOF00LqQ2wgjq+e94jIgTEqYY
aY+yV5puFBKEWwe7tuiYNbZTyKaTxUG9J9iBTLrek/i7vLczclcpTuj4CiaksrXdNvcjZz3nk44r
mJXpIhxTRzFEAPRie2di5aLsnJ3ZqZVa9N9hU2NkWZFKLl3ttS5AXYWVYG1TJQp8c8CuEom/4qQP
Ii+/Ml/P4wXzi6uqSZmIDleXIdCSfEGTzJFbiX5RZbrOQ0AbgFQUJ0vU/28QeJJEcmtPVw6avDKj
a1tg1pxS4P+WwFYFpR0Fsd8VszqphPBo0TCNWhmRGss5AHSEeyFcbptSostwB+OYEBrKuO22P50k
VMPibIG7VVkRGQFwscxnbGbHwKiXL4c51dywZu3Mis5mC7Av7/1yAPN9SKP3lWOiqz/jh9+qDKf9
pQ/EkvpRoegMbUiJ4KWx1vI8KlEy3TyMFtWYtibpj6HeHkbLF1xX9QFKcgrDBu8RncUwTnuomIRr
foczz00t7gUpNFQ8hbER/3b50BxIL1sx2Wn0p+b4XxPlodgsQ9EXWJ90BbhXFfZsq0Cqln12kbxo
qI+09OwyJyCD7E7BKmemGnScx1xv/deZHhV0D8nE5LIf/YlLDGM+N+yXnRbr2EWN/GGnoWK6cLg4
rkZn5GLHwy6+U+u2ZLChGZsp9eGFPetOeTXkJwta45/JX3EQia7Ki+5LwlnjeyF9t1ajGaw1hQxE
tTasQt1VRXHU53a//YrfBGBNDc0TpsAk0f8HnvAHmUuStwwn2CmIYXJFNqJHdC7gqFO22xJZTVm/
2PBrNAmgSoIaapt6uzDXA2JWEpa4aOHKUxPIIz4TofUou/rWfIQEgnWwhJWtmGNBSKQuryPq3ahx
trrdOMJzN5vPDso/g77CopyewYimuUsBIvwXcMflPhZb0LsSsiCLQUq0x7y6FxZvj3PLQGSjTgcv
rMdui1L5kdUEGpzY1HEqIDkXBpxCXYn8UC2Pqlq/KPB50DW8y7wvWMFJ2DnKw1+968SfGN3pI4gF
Xtv+QLxyNkfbwQDoDP9zUPogslZSZbh9N/2luU88Xr6m9HDLAGnOscGxeTTBonIxfXac1Kf4ac0I
oOm9GnKE/wXpIzC8auLdyYbvIEcddoCXrFCie8qK035q0730OFaQvFdhitPDfJ4JGLXQiZIjRa1J
Y6uNJbhUDroiAqOALWNxS5a1hfUp/8w7Rxov3piHllrK5/HgL7ha1/WsknOGjX5ZpAr31QtE2jEj
F25FMUK2AxzJ+WvNuYmGjLBLdmTiHhzMia5IaiCSmOYb244mRuxV9x3Kf4dgS6azzl1e9zJtaXga
4c4lEFtG2avnbH9iC7KDjbj+1nNVBWjtR05LUkq7BVxjKM6zVYDfLNZvb1elfJ3puhOs9yWWPpDa
qsqkRT3KZJcy0Anffesz9RRa7dFHzHFV7rYRbK4S8jCqJ5CrFr6uYjHdKXNFuF1PrRTj+t4u007d
IcUVkuucdG5ECb51K7aQr7BA6Xt88uquTE0/4+wrbnuvYRs6OlFkRpFoD+JoeLYjtGw16P3e7b0I
oYyXheV/Y0r6MIF9AefHiE+oR1pUrww6llZGUFZMZnrKGIH2AVwgJ/ALC4BgWUZ1hMTAsIDajTRA
0JnY8kC3J5yFAMZ4gkLrvaCRY27ZY3xvjbBWKY7D8tIB7cQRPRCfIJsLKdBr3n3LXrbdCE+oga/U
yShLM5dMCAgBH0n/T+iUYB61dGX7rQj0mKzftMrrQvng4yAyORAmj2JhqLDhYVrYY8grKIrkPbAY
qdunW11E/2+pWjiS1cCi7bif0VswlBcA34ggLZqEIgM97D2oOJyDpl11nG3S0g7CZd/U13X0ae3f
RE1pgosXLOvC3g18gDmmCxeUd2vUE0mkn1AnYA/+bnK9WcPkkZwqS9ZQdisLQyJW4YpkDI0NEyvv
JZUlzR8VWOk01xgHZ7PKvsnVU8v4gRpeyJb9bJAUYfjw6Y5HRGBKl9adwSF6C2JRKgapkpF0Egy8
jaKjy6hWwxyDZgHinhISAzxXuMuo5E9zcMzBzcKs+9y0sSb67GEL2jZrmdDhw15fUp3nWWTDqCaX
xtPOZm1yi+430TJDq6ymHC8HwA18fxziBOKOZfmqbf9XxFNlQRM4HRXao7v9neyoKjJCHOCvtwMH
qZAX1x2DezX85s6fLOX8/XdzH5t4dX7zUiZVaNsKuH2sIeFlb7RtN7/EX2PNEL2VZQ+QOwm7Btt3
EsrY3tt9E5hwkI07cEWVhABOUhi6gqLxah+cWUp5zVmKtQTmcsZcNrygdyH4oaZen7ROh8t3n1O3
MtwZKkaasYxn33TNrV1KytvFlF/k3IbBYhe/Pqk/L/5pkBj1QAOsZV/g1Hteuh5FNL1tSGVekpL2
2We/yKIbqdPS3VP6BnhfWRYQf65rNLajIhLZEtncViuQ1dWVvIcuCbPl8wO8KZ6jlbXfCRg4HHpi
IgYdf6M6+dySyvzXj3xlKngwX7ZAgijQM6GkWxas/Ap5z1+1SP04MCBdC9lkYRe1ooIAsQ0uGzJY
+iFJGrhrF+jbzh0d+zlHD3wzxvC+35WbwTFKTQj13EnsWaOPr3nq4JBjZpVWp79j4v8vLu90/Rxi
+yjCLNGtJ4t0WX+80WRCpWMFDg9nFGmLZeDlEXVk4iGy4+ScA/WaSnGRjkmal59IPrxF/j3b64ZK
5uYO+7Odnslt3velso+W6QsZma/wn6IAbh5eot4/mxE8xAOVNmGpx6GyU6QlvBWhvggY6T5JP7nP
J2naCE8LOkrMsNFRxiTf5rn33lJvLTpUQdYQpb5xY3H0RxBXqRktHzjTbOyRGzyfeE0MBp/SxRXF
WPqMt2gR0VRsbm5cuWMTfkf52vLYXusX00JS/ObzDthNHpfu8wBzXuxnGFRSw70h0TKn1rM+kDCK
LE9dvxzRvYivaPg45BaIOQQrXZVf/9Uk3DlIN3cSmKjH1RUPhbAtavoTpINPnNX6jkLVoN+Yusi8
I3aDkNLX19RZlmXuLhujWf5ArFZ1TsBTJq1j1KVF0uaFIKRG+mMd6A/v3usd47kp4GzyXbGXwIRm
fYrUN0IIO9x35fdUy+refuebry+Qh1TVzwfAL0/fq3FTuXfPtbU42TEUXBDkraLKym6hD3fqZcEf
hFL6g9zdHsnV1vAV3579pnlfMwujL/Pwlg6FsQHYLUKP98HME3AK6TmSRYXIXY1nx6N3W65HDuFc
VwjSrqLJ9gckqnztXIzGK+7szUZmtDHxL/G6anLyC8LWSs6lr8sNr7JPfI4ZFDemCtGmFErBrHnf
8ySIKykZXgcIJC/vPjKkEDRoA+Cn3L4TRuYJpy/2Zv4utiXIf24tIx7FN6/yFdrHTsJNWhuhGywc
TTnYkk+wXcrWGAFBeXZ0I+IimBKR9Op7hKJx1GydHMiVjsgYUAG4ljS+RepzZBiZnwZ6o9UZa/pS
Ns5GsQ/cYHcyBwZtn/P6w8W3Vrpr+9z0ZegKbNqRlTJag237Z7DL1crHaPbd/WDh/61xHP+qXEya
Ui0WzopsQmivviM5pnK1rwpjT+iMNStAPUs2Paf++6CDxFvfJ09fLsIFy5N6XBa6xqHq6ELgYe6S
zpvsOne0NPbM8xQVkOQzZQWvsa1/wOKdXBe2HEPXWKKJdm0ikqeRJioXaSUhYAEexn+86Q+cX1xA
8K4nmOqy08jRlam1R1396S8hnMTDmuDWDjH1mhyICHPb/R7lvks36MqMnu89YrdM+W2ap7/sUHkP
DPpceUCpp1TfGqHvN2MxtqNt8AVCEJUSg6I3eByDcC7rYlqdOzkUuKkZUBdKuDTbl/9eqGhIxMpu
U/IQiyTY7TP4tcQsjibG5OXu+y9y5RajPx1+yZYCsczNT+uFxsIByYzoSfQ/Ocv8uF9JndifH6YU
jBrqG2ePFcdt0SjTX84Cvj0mBcaNBa4QVLCRT82oM9wvk8+kq7JHAZNekIaYoIRWD5s1xZ+3NJVN
9NkEST0oC8/Oe5E5NHTzdIoQbVKPYzSKK7s9icWj0Z5ceepD/EhNx6LBdjUMfVgxNLaQoWtBH6c6
JGU0EwXGaJ6E2zOD8bEZbzi8ZIh1En0CpqbNIfYkjEXF+BMOHNa7nUAa6F+cuPgBnL/Pa4bpbvKF
BLtZCyJ7Fs52xC2ShsHaH3WY12qnLpDoYVUthNgzxqGtf08NRxKIOOyHh/or00/lRomOnf+SotVm
yGmLQYGV4PJSmSaCMec9PvuF9CgiYPaCSUxew7VB0A187QVQMCrGyZxsrBReSRFmLL75ENHbyjSz
XfcZ7DdXmZM9Mjr9El9n+VEdOGzl7+/qQUzrFACsDcvknDkFhlXtXxjY2FEE4H00ElgJ/TFl0h4y
iejXGkxD/F2MFh3pNRL2wgoQI+PfCFz+keaKts4NTMbm+eoi3/VQQLEsSlP8VYonPdEMTnfjPXNl
2uLc4FKBzpDFzgiZrMCyxhM9K53RoKmwaalN1uIGdQEPmy/03BJYLVLzve2JNiu3LrmJP+RjAige
oCqsNcLzePDR62CCiGa3Wkrhndi5uXLQ3HY5cEPR8KJZdYVxIfv9YGHUyq7LIw5OqvSP3IYEYoDU
4pThPx10BIJHZjTKr55C23YGdnMFkss/VXBvXGdXXrvnXX4fReu8Fw1lkO1F+01QEuciOJm4Jt/J
Phs/WAZox5FoXPx4eapx5+KIn2prhntmLB1jqrl9IDASJAQHXY7neLY17apIOgTmoJk+/t5U/Kk4
DP6Kr1xeHscks73PpQnbdiEMNx34n/7xgw+tDpulNnIhPFHWcY3/tMZ0LJZmv73Y70f/NJdFuCeS
KceqN4mSBPItgAZ9dvrqxYhR34BKQpToA3rVjhMjDSrYDpTpa0kJHoYOA3XCmYcFoP2HXxtLFLbt
LsYH/0bbPS3xHqUVFUewl8SB5BZ4W06t5det9b0KtloCU2PKqmdwV21dpMzZWmZVNH0qCGhVYK2a
ENd0IvXNEUdpL/rfkFm2MOhSsEySkPK4ArBg0ZjQYyOwTTZFARKbY/cqLckB7EqzFU9YkDrO9gEi
YRCxbePnt0tjaXGt5crYjyCQCmEM8jZpSetZVImYCFKIrFY7Hr7BIKjonkD7UhMTmyjRP8huxn7l
vQ7+kMccSWPUowBaCzoKoT8FQcauy1vwIT1bFN7Yq0M9QkPmyAWgDGG1LlrHUdp/CwMS3q0+oc2w
Np3Uev/HmqAf1v/Src/AYzthXZp5Y3OZJQXpVoSWWdWot7nQlRPdAUsbg0jvSVLxfiTMM8zL3hxS
ZRMKo+1HyKQy2hj52fTD+advWUQB5eVKrre43KPVMSpwKCBcaK/d8vIwG+ggch5oe7ZRSNsarykC
YDNBBX30Y/MfdGzZ3ovd2NZgjGRFpg93cxboA0sLQphrRST28DhEC39bUs8lTSkX3rHeQXskrB+Z
EOQsYGq9rZni6GvH34A/QdIWnvTl++PyWwwgChdXOz8jiHEjQbEM4gLumaewqgD3fCp+gbXLUHzj
CSBhhR1Kh3LGn3VPYIzAsoUnEjQ08mB+FNGItYYTVGrGVb1NrHmtQpQ94gFA2kvatJnO2NAht5rd
f51Ckc9aujS5CqRSGLqJXkJj0nrx3KLF+hYtlh8wteqfv0FIKimcSuqavtMN8tafQqnsCNREopW8
ugrB3BHjBy3QybN04f62LqJsIdc8OdVcpc/IIKo/TtxZQnGaYAA3BNBJJ4z/4OFXx6Iw0NIU+Ho7
KmieMOTpa9q0lu+QFtJd6h77fag5n0g3GTe9rWmH8bJD1vf7IA0LOWYB8aCQRV5JjIab3djMOMib
GkQWj61ayWzgS1Ru0S0lpUbbOkqYRvdi/kr5Nv0nYYhrQKVGla2PiHog4jlHgHtkaoqM6kCxGGUn
b8+4reBuy9qn8WXlnoRD91JekHAcpsfs6mBPN+LUTLclRv2SBzmMitPHLUGuMjZ6jiKVD5cZsnP5
Ac4+1mzM9kT01l04vaEKn/4BCV8FT32L8AfQ42f0w27mBUzhQHViQfP/ioZj8OeQKvj4ockDy4mT
NsDcVCQnWWafHvnynAIUxhXlsnFUSvcabCyWEncS7Lz3RNVT6PeMyvix+yNM/ceh4JeWn4TD+Ogj
dlfSQAmPTjfvzslfyA1S0czMaT3+0WwLzICORykqL0kA/18IGq+yL6RhKWsKhRCbxIaX+fQzpyR7
M41l6UT6HtB5MMXc6gNw6xHM5IfEiruvm8YbpVTk0TGTEsO7UBw00T13qujV0DMK09ckTBJdyzN2
B+0inenU+0W86MGmSvwPs55dBByjNQTmONOqdZv0Q1VF6uL3Ka6lpuIRe3FFDkpfbq+KKgvtKwu7
h+lVcQ+vi88eIlvcT3pPnqdT7CnzkCAAhVPF91+qn57SRqerDZaQg/U++lg1VD5v4aHaGXGUUR5N
WZ69TbKwjpIAC3fUbQ+2BRCRBAoSSXfAtvDF9cejSpZzuH3loPyJH2tzmoUjCxUhORH2p0xQ5cxS
/8WdU//iP6clUBYMF1gSBQTeVavxbuNbNMhvYZHnLCnisNhrkCVZIGgRIVCztkDN4MRboscbmokX
Obq7tjn6307Lhtz9WN24/hs+XQ7PXktaXKYfOrle34ShOYZW6uWhcsgDWX3A+Z+Q+XqR/ENk8lny
3QcnJRn3Y5xUBTitCxZHzr791iY90KOtChZvM9F5j3G9sqxTJorDtUCd0kELojZttDeoRouNW0qJ
Ls2a6p0qXMvF5xueYgabJrS+0OQZ8WlVphnRgK0tHPv6TFkDFcD7jW1gfJdEHrYxjFW1bXTQHPLa
yp0vstBA7gf6O1WvVyVKzkohKmu3Bz+edJ69/tGCvI7J2y+q0Daex5pT64cTsv/dPvAFu8xlQIU9
XDTaBzHClgtEImn3NNfC++st0XraKWXfPh9ytyQX099ZPDq5HMXgKdJCnQUpUSP4vjSViv/8tywy
Xi4V6LK0KcwC5+xCcbbWJuXKMf+Hiiu4chdAEiknxrt7RoD+G5i4mqgK9hlQ3DKx8DigiSabH6yF
4kAbfpKKGKAsYV+RgivAsK1sKFK+ViN8VH0uN/UbIfDvdrsbl7XcEGP41gON1y+iTR9DkllXyFq+
9fSE/QEPbb9z+NgLPzScT6f3O0QRlaOK1x8wuCDK1nZrn+wYrFmrSRt5V1vVrBVEphnER4eAmh1O
AdmV+K0JLtKs7yIFUV8Zh4PJLQe6x+QJ+SoKaPPLLKgqf6SD+KK5OCkVawA8Tquj++F/rZktEd/S
ESGDUt7l8zPlJasWv+ggM0D2v6adt5IgRhMkMg9oi3kBhqgyw/GzIzWEflc9xzNdptrz4nViFZQb
8EfBXR/CdOkXwEnY4oPenbzPN2V3A9jXJU3xEPceJEQu7aSWlL0x4Gbp1ZkJPu9XUspLlRW+ci2M
rkftR66hIo0eclLhkiFLmGM2BlOFw0711UTnFjXJoG6i+64UiBoNiGjm/irU2xxZMVmjYTBb4CWE
YYKiOx2898CEdam5VL7Ux6vtAhAVL1+Y2Z0GsV7axZP8RD1cFbC9thVQaooFV1KY36zBEPgXm5Ot
TqgZZlaCMEaBSpDP2j61wHVhIzzGVJpirXuiTFBAkREv3MOr0vaFvq5b9o4GxywLm6LRk+XNteYo
rvBA3FiNfqkQJAprnv8w7Q7q3dGgDjKNgm+iZZgtxRoc11LHljo182SYb2vhDIQreAgcGDH9/KvZ
mdjV6fbh8/vrMRknL5ochT2pD8WYqrvWyS0JkiS/0dLrFkPiIJ+zvM2vDcnsSqby+sbaz6nEFN7v
p6RMdXICKtihLMYUb1Zz9a818RBRCBY8kEg12vjtTZ4LVQQFrPzO+aaZ9weVYUFGwOAt352EnNt8
hAEEZKT8yCVrflsR1Bz240CkgrAv0xWxBpLVQhHeriwQrXO87H+j44MZq716ZqEM10L6gvhoma7D
PFQuhc9lo3CSGwZb5K8/1hT9+4e6akxV4trgqnR0HiAt4s7UVGf8nRPk2HtbhAufBXLUXnLzQNiG
uMwDrrcS84/Gzncg19fL9zWd508hqL+Da/eS6KANU7AQa0/wPVuVUg7aXSomKVWHIwwA29+EhEz6
uk9oPMRFdglv3CX8SP9P2u+VSUYJSUwn6uYH6iFrwRQfCNtO8hbzkvsb42kGKHZopMlv4giGOv8G
emflq3vplt9ZfdDt3YXXPk8MM7oY3TtQ3yv1H5nhjhZ+qtvJcst9vK+feexck96MbU+Y1rRxw48+
cI7Oyb+jxkxtC6dModghuvxWr/nKOQJSJFPjBtZnm8HqTLUiz+fHSz2OjAIDTTvhVz+XYlqrDOsr
viD7BaboOkprBfjsDH7sSX6m7srkpWV4zSY2O08M6UqRufl2pk8P5jYZLE9BlxPmTK3PsDnl31+x
an9sE2cQt8N0fvYo1go1eb7CQedVHFgJyWzwQxXszPJGVGu5Y+yZGG5ZYF4KMSNcSmGDdTT3n+9i
s4KAFx1triYfruxVVU7unYJrpLXRJjFVwamO0iypvJn4Y5L6RwzQEHYaYY6ofGop+0uDGUtvF3hY
/T6r+12/6/4V8cwcrXoBtNxx+9Wqu4SWVFiTqSPxHRRwl+VAepLLQbP0KyFfAsWzeYIi2NRKaLYu
T307UnG3QNKsnzC3NEi6E2LVHHCcJ4HAaPYbVwJ4JleyN8kwXmKIcUcWLjctb0RhgUEQVkrLp+4v
RpDVAfPJRiQfeoDlmqzbPsJIzd1wdthsYwT1QdVRYTu7gjpfBTnL/0qtzVGfuxU1OzK+RLP00sZi
pXDukSNlvGRF8zn8T7CtD9uyfwjlh0iK8xM9Oagmb524IxU9Wiqfq0hUVjwcYSJWX6loUdCSg2ch
0d57OK9rIVED8MhF9U5qz8lproBtxOJx72j0tnBGTXYIshmDesWwtnoyQPMD4g90bLsWfm+AKqu1
0x9Gtgb8sPxLjdbospSJlRlnEFSZZZxVdFo4PeQkd0Bb7nbGPd5TmP/2/fAwTkv51q64/P9vcIIu
+DLQ4SfVdNMkirP0xp26w/dzIs5nzy+SWh6LeZ12Az9jXHTnp2N0n5Q+FWWShegqlLTk0mKC5XRI
VHQVl5WE4r5H88qfnbXvn6xZP+OEs7tXtSN5UdvoaJbZnftXRUypcd7n/aW/Ghve7LdK4+bmsxIh
qatk9HVDzpxS085EF8DPwao60HQND5BZfOA7cyFODwTr3aMnaYoiQi6c8P97zMQ3KhHel9VI8jo3
BK0pKZ04NoKyPZwLhYYIBzZPy0nmPfVUj/4OA1CFAIaHSOuJJePyP4m61O2af+0GVrBJl+FDG3qe
nEgB/+qjqKu9tMpZPvZmXPb66ysGfI26VlITEbLSB//x7/Y+5hXX6XKUPIKepVTVpzUDKU5kaERr
s+cPBaGUk7GTrRdtT8Sd2A5El8UcAqZ1yb/MlXbLgQzvLJm/XhXE7P/jVR9gJZz+jJ1rx/qstDCm
LQ/4+vwUjDo/V+6YkKGfu6lL8gVBw62AHf4FzDWg57MBLJWT9qg7IpMiAexiDQmhSficT91xJTiW
AEUCzQZfJxl2en/1XrZeRZOqph7gNdYtFVCzVN8sxPfAt454cohnHEAL+z10SUdXm/Lbf86xV9aH
QOdiucyBRWIUmONecnoD0/zKOT5vB0Xzd/IdeQ85GFWlVN6rGHKDzn92mVKiSbqjlHNjZT3XGtWP
O1muVL1BqRS7zaGqzQSLnniiEXUcq/kfaG1X2VrLglsgW4wTDCJ3TCfbH60X0dgDiVeD+agikCcf
IiskfoAa0caWt781q63RicCXNXnlkZwMlXNzaI6UnzRfwHYLZ0sgGjv7q0sPS0ZX53KwNLPPhhpd
I/WFXiqVlfabfck+q58OUk8il6fmiwsVENvPKwLPRuIUWP5TL1D6HtEV4rcQ33JtfCFOlMRu9c0I
ygdsvV8m7OOLtkjiJOWYA+heq8blr1Qb4o3Hzg6BwP+7RHoan69tqv2KVxjyao8gmCpBg6gkLYWA
q24c+IX0ZMCUyqTK0R5b0iEEBE2iIuR+WcHa9BZpMHvEPluLop/rFfBGvqOV5kejG69ioTSbtbF1
SWrC0ruaVQSg//mXAL72C2puCjdwJ4qaB4FKrhyqmuAntszOc+xLihi430d6it42ibucpukngpXa
m4VL7iZj0mVsu1B/rfCWJTvgSYofpOTEsuV2wqlaNt5WRhGk/p4ywn0HCdx8qr8nThmLfKgokZxq
s2jGhgIEUTay3GB4CRJ+9eGfNcsNO+bGBIrEpNRyYiDuMon5OdYOXy0NGuqW8ehZ1aBOLG4BExlK
REy2/sdgfOuBzRMEUmsnZd+YMqcILzNlrn9hrwibbvHWbOvDi4jckwgl3cOHfamatgdXPy9yVu9K
l0Hb/YTeA8lUX6ZS+A8K6d4XnmnhhThsYtjljYhUwvstcgEoR8spNj/mXktI0T/lcf8aQGbZ1QXX
fcP0wasi3FP/tzAYY6f3+2O+/d4r6dOoJM+tI/mkcLwdyniU6Q17N8XXSGg4udlHJfeEPn+Cb0va
GyXikI717mmHxd+nHtIMmwe1eXY2EnWuhh0H8prBayNSAmVdjhPzKZyCjCYAH5dvrfW+ueG34Wrt
sDypxLmjo/q8T8dHNxCCTEw8ohmm+ngadwF/TW7pN7ZXr/5Tj6yG9RIFA42amc3DNgYnE05TQ5Jn
HR6epwe3m0BVXUfw/AP5d74QVDqbkU8nqXcdNygIRop7CcVTQ0hmrolQf+z4BqxVWhQ9FhPJfdjv
6+obTLkkj/xkiBc4AdblE/OkBzjRIdcHSAVdqVPYLYI8mADG8VHGjjFwf1C1WkNFp7n5tJdV+2yE
h0bgvSeDn6Aa0OyvT8S7MdVizA2dOYUFd1J1i9k4bX5SPaKvGPEQxJJzcp319lCCsxFlfqdsbiA7
yQFE5Vf4kGN8tO+tCbzd6WKNmMh9bYz2MlrZeE8DvUYdIsPhLTE5IIOE6lBgCw5csJ14rMnC8e4n
c2Qqao+ay8vQWzzdbQ8XWlO5KyBu4g1fkuApsEa+UgRHDXQjLf9FXSKL/UqKrlk6ptxo/++O2XAH
3/sZQw/w6t/v9p5wTDDcJjokgPq9p+EP43CgFFqnuHSl746HnW1pef9QXjAUerjUJY2U9MtEdp0H
fqxTVLXr3tf2OPURzbLR8dr+ex9yuO872XzVzgLxFsf0scanXXR35ad+1fanCe7VJAdIwcUtlzB1
AUQUw8fNTEedriVrPyRiJkkjiifZuv7EsLe+ecuLo0hykzdzlOJBbqXvMWfjxyGANH/YTgTD7kIK
s5qAtcKd1m6GvoykDibBnnG9xgnRjLo5d9VB58o/vlwgOIHB4RisRrpIB6L3El28lyNBeR/ftLaF
nZmRBhqTfXBi4wM+VN1X8i7N/WaYoT/W2JcuPAcToQr3NVVpXoul1HpNT9yjroaWHoUkqPapN88m
fEnBRxZxclWFX0cLUkSIUExD2arknxoLjzJ44U/z6yMg1a8tLGhi55N6LZBfEzL/uQJHMg99pzw2
uoMySfb1QNDWVS01nwaW4hghCKwk1iTToeGERpCWOWla8ozHo07nvDfTSpSN0Gwv4nAHVkPiPIhG
B0NFipTP7kfjgIM+Z6a1weUrmNEtKzY0UrOwdVm2lJ10jIvPwHQbRMNRN2cqsPt3F5sGSe82WIJj
dejoJaOGvGhXoBenPgYTBSKNNpZGIePY9mK5Zy8NOfAuEz1VdgCJRNAduHjbPUffpNsNUIiT/pa3
wtz6q6/BxZKI4EohuJuoRGvS9C+1O0B5kF7CvNZ1uI0d/hITP2a4/vsKo+ilpSOG3lahPUZrBITA
yKDgItbafuBM2A7kMvVU6ODEcaBoigbQhmm/PHy8bpTzrXk8RrbsNHrcS4q4I1jDupSClMskzdfE
1V5aaJb0rA7EJb8CzzaZ+tkHO47HiVw6hDmslr08SQ/khrYx/AKhlh/0/DFOoV9PiqCSEhVK6fvE
c/Kh/D9HcxBsMeZFWjQE4UDrhrzrzqTs7wPplfSaI8wJYrtqrkswfeJl6reDl/QyCULsKav45GAl
FKcdMW3bkWQHCiwFz4lMDS7sNL41yMt4owCSOShBNR1k1SegJxj+UT9O7ljOKp2UR13g5plR8qln
2nAmmAvOm5MIPYnw+XEJ123zogE92fRGpvDgFaC6XJfMb5YAU3AeWH23xHCGulB4j8/jbyDiiYXK
qLkggYI2EX9tXPYBMnPNowfsbjDezH3zfLdDHpBROC44Jzc+uepXVJRJP8xM8Og9IpGMVZkA54eX
UxaF4kvxHN7yMrVUWIkdh+ErAm95zvWlQTjweRywHWO5JhDbnto9VMMwYfzu52H8Fk+mIYDUq5oZ
u9geDvVnPNj0PnaUAq4HtijEmMWF0fM+FMS9yXuaFMb8C1Ai/0oNJT3yfU0dQZ0XL5/g/hq1a5J1
BD1Qm83lL50TnBJVngJU5ILJhoxKcnS8+m1rFqemuQEDOlgRAkEorDZzjMtDzg0GRnzTt8ndCa7I
HAa8K7stytIUP5Uu5n/mf8g80VsCsZcRriwWDPm+I7SYB58YtfkyTpgh5l50JmY19JGqSvVaOrMT
3XUTw37VJ48yavoiLXUNHssrDPFWxbqoND2ctpNp8rYElxDEKIxfjYT7omLHHEps0CszRzMrcgWI
jwbs1VsitaFlpncALAhIBbNpiaFnDFyeoHqMte+Ji+0AUhj52s+83I+NNvhtNedi8vPAj4LQqG7a
JsfVzehDZsTKFUsVpNT2m+CdLpz4j6T7lDd/LyID86K8eI+OTOEV/CZxM+VxFudbqfiE0+bYksyP
R/eJL2+Egi7m+olr2Dws8iOUK5evhcYt4KXKKfOeavoh6nC66BndTWPAnoAAqQBBuoY0pzqy/kV1
XIARX/ZzM2/5r+d+ULUdDhSPfGIvA4prdm2TdaJW1D23cB/Hgv6iNgJQ3nQquebRkoiuY44XwGZI
Ug66o/VivHharEdYJrexVwQn/AS+8mgDn6ZnJLeaxALhrN4nVV9EMCvP6Ptu0OraATKW9qcXY8vc
Af5eMJ7T85JKZ5al5FJtXizMumrSLeMgKekKrod+cEPKo7P7PyQE8kVfnbScZubylGd0wXoU4GZ7
L6vquWvFq+fMIYvbeCNFeuTS2YF4y8CnB9QOS0SisjUoqRsbXAad17mfxafMqhqGd4VuSuSGY7eF
AuxpXgGTXajg5kd+Bc14Lf7/p1Bwp6midZQwz6gIhy+qrAV6wnpKGea6xcj+SZ9YpUrskthdw4TG
iXBuCaZ5GsXmcMxvcHk9GqI7vd8pG8mo9t9bML/znQUomLhi56zI9Axt/hzGsABbpNMmmvS1oh90
Ig6fGXWSZf6hGYpem2dIhIzQBiv9Drb3Enctkt3/6TGIwkeD0DOUFExi/ogfTWjRK7oj7NlJVs4J
90MlKxkjS0kmX0lPt4jndaUtIwpjjgLitsI51VKfHKBYf43mtVFN6Gt18AzbQf7vfTt29Oe6k+cK
THyad3sER/EjRL/edjfg+yD6YNnuk0oj0wzmPCykwj24wm4hLclyswXovCXCXaXzHS578kj+Ntz/
l7gPBxy6NrdMII6nmISbInY0LmLo/0iz8ECW0Z/05+iTnTF3ikek2nIaNucLD9uPLdxx27HrOKq1
DDJl+uKyjOUwOrI5CW1tCxo/CKp8U3VCa+Xk6UzAnm8G6lIvoAHhhqqL0pRDd2gLCKxgTvx4l5T/
t9FfR3arme6xxJvozu53wHqoT3Zc03Bip4U8QH6ZyECbY44DmjN22tpYxfe0IZ8/zcwQAf7bq4B4
gG5//T4tf2FQ5U3k44M4E1GUzbM8fh9ftQESnHLr8wE1mfNLHbVJeJ7yhdgWvSERUmcqhWWMHuZR
ZFPHo15jjwCH+4bwIQZ8u2ILN96WF8pxY0/miPN2F0kCl8N1ILWpCwF7xNTipfA8DO7ngcqOOi81
2w5QSvcjL3bWMR0bWMhO92Mldwg9zjLbfdknDtJKTNHU2a6wVcF/7+XUd98zuG+7tQE30ZX05xyn
JJs7AZe1LWTUw8l+Ai+FYyDc8oCP2w3QkNuhGoLRWASnBFT2Q8y9lb9G3bauz6QScYS9Demss2Tg
7At6PcvLPEcvFvWCE7cwabuke1OUoF9Xy3NeOpwACGrKhhV2wDAiv3n7egv9RL+gMh15jACOYD7E
swe/bCaXzIS0J5Kt9G1/QCfefr0EY1jKMrPa2XXOIDCqUf9464Qc/XcYuLViunhAu/ckaqRRvwa2
/pVSacdiKEdmqi4Vv0QXsNTXhamcL8p1f+smAYZbVnGupy2KXNhO7qsuzoe3aqrA5Tgb/+gr9nmp
heX1HX8gavpPWw3PhdiT+0T2lXRDk2UhPEhT1YN70ScqH/kLMvmeZHOjHoOB2mxrQpEP1BRihLyl
HbaAHOomCaPP7UlcAVwWmbGWZzbdcnzIw9XwO0uq/zUBOnfpkHTY/Y1I8NVB+4ZnBcrYwqtt/9/m
5Ok/rEMhEgkJf0xfmOfchKUHdd3Gmr9ATUSgFLF6RN+ADd8amiV/Y9n3GWr04QA52cG739IQGfHW
5orOk4lNqLqZiEkd1q62T46Ohx5TLQnOLsyI3Kg1AAr173syTyD/RRkpc4ZwGjhKNkM6MpFJ5HP1
3qs0szh4S96aDOR9umUQV622yB2OK0665IyMYEXzB8Jf1CXFg8kOBNAqRkSc1WZy/ibjpNhVP3R6
TI3E0XhFWLQGLLSUFgeJyPFQS9jeU2sEfJL+AmFbYy+NzVJOMZgek/Eisl8Snq6+7ZgQEF1vRpHC
iQhCU8EJXojKBCSKe9+nAYlHZMVLzugT6zJjqEqthUURyr5ryLDYiYYdSquBP8HV4KUpfLr01+MR
1PxlyUlHpe6LnCyA1B/DYN2UDUyh6nW4fbBIvxkhiOxmoH97XJB/3c2JLz3WQA+XELBaxMoXftd5
JuhLXEI/iTNdhwKd1DQbbAa6NrK5bDSXh7FNFrhUmXCwqCP0/IFq2dT9EKKPw9YHj/tUl5eAkCrX
kDuk59GVRkc9AwvfBKZASbwshFFDRCX9luv5MKb4lCgW9orwhHY6uq4M2ufdfxFK0iaYByjOgmxH
tqfjJ8HSqBoDO720XRTkAo18ZiLIZfYGD+a93T2Og7INrsLCsfoLAOugsSK3gaJkViAgUmAvUkHk
/8TdWxlGZ6CPfYO5GcXrJj62k9ew62BzOPKL7N3LrgMGJ2Bu92JA7J3rdQ1FFSSoZs/j6FwVVXMx
GffbODGsE54+f5tZ6XJotK63eW1b/DFdP9FUrDi9lFshNhak7V07iy53h9dlawDnJdodbCi7zeUR
F/X1C9CoIMoLkn54+Z1YqST7lPaQDSFMLOiEvUul0wyzbmmpeO16uMUssEQcM9JjKdEKfCWbG7vX
dZiWY3qIXcTIgiMSv7/w/FA0LmJMSuetZ6wQ2uGKx4KNg6Xk4unzaA3MqkmSeA08FJO2+1FDNkxM
f/yTJVd6ZuhgTHU71pH0Or5iucbHmA39oRsNNJKAfNcXXPgXRG7cyV59NqEN1E9HLoZXPSLOug9y
ZgtGAGBnNBpNQyCdu/2/o7HrqJfu9ybf9pVZAolEf7Kf9Yrqeji031pOSmGsqjbBR+We/ehPTMeu
WGCYhdzgt+WjpJgQ0hnRHgZrsr3TM6ipAMAq4LfXrmYRFgOL+MOAhI1OIbzT8EbPtkP4HQ7MWXl3
r0SmDS/tbfmPIO5RZRlNxWkbOl627OT6H8nHFogbcrY4gmCo9N1oPlgrSZVzRusqPAGOF+Y9sFUC
/bDB+EWquFPJLBnkREsf9o12Z/bv1CRHDdXvdX+wM2ztv3HiI0girftIL11oLzUc2DkPvxILqCns
GFC7Nq17jQhWT3wjla5fhQ3Y3ezx6xDSNJZc2VIfLzExx2SdgwvIxgHAc78791Tx3H6fhBFy/Yvc
Jb0ShlSl8HFrLq7T5Alzbj/LXEtSqa1hRKhBz+pv55prJi8bNWQWVCPC4smuuA0nXMWY4r8jpiwx
YpTaiI3CQnhuhbua9e6wwhjXwzj898PduQDneCmNa1d5UJZj0ZZF0HiqdHkSXOVfe2sBLRuKrSQX
+7hSPvpbkgiSRfGjcc72K8Tma0ZAVpCAHe9JHFZFWNMZ0HrxyFWvh6T2oTfcffs+//VGdbXDSj0i
PPtWiQBtkQ3nfdQ410cVExjAzALC5GQy4r6NxmTmV3SnCzF/pnVGv7aUZiAE8T/xgPICUeoM22gF
jjl0ikquCdNVILGsnjElQVO6ay1dOufX9OjXnpBlvkgPmLew3fK+diuGCFoTYAj/eyV5cu8T1/M8
TW2oIzeacHm1d+4TGoyk3BkPytDO0xKH/odOekL2ISVHLA/474YpsUPXB5x6Q6/hcxwxTinMFgrV
GfP8XaN42pkzPHQ4A8AnA8L7gLObRIppXP0ORQp2ACEkG4KN6KlHg66M3P7r7x+SJYWuJekJWcFU
/+OPhFbCNjGuYi8d0nzXjG7dsjLe3ZYgDnWq4swKx5CocOo9MKoXHrfvnKbME5WuspGZQFO/jR7Q
Db/UzA1calnGvHSC+ZkVYbvEiPU6foUgo8v+K93eOki/aKPDamYIZhSPImxuPz/MdtUZPtV7FVwe
/H7JSord+3tlxpIE0NZ7A1e7vnuvZZmKBRHl5qrmS7XCaiaJLzIlQ78Jz8PVWfPuNCCLp01jXdpb
t+DBTuM/VhRcxX9zcR5553FfoCdDjsFASU3F1Fj9uvlMqzRJhgKk0txsiWMpA3ijl98csWUzyJiY
Bgd2vgeHhsIs7tgxToJmHmSMabziHeZCFOvcbhMtAAIhn7ZvDhWCpv514Dh7Ijd793tiRQXqAvLl
pLyKQAunPwhXkrVND/+OehMqQl02NtRJ4PeJTQIEV8ZaDAC9WriCQjp1mLQQHOIXQQAsMx1UCLwJ
jXbe+sCmGULrwb7omZaCHpd2yZ/4Gne1FT1e1xe+lpbsKyZch/xCRa57/9ClHYvSIxTyUBV76msZ
NNZ+7+fdW9K/76ZdXBstK2uxSlzjfZ+vSHvvfbOyTXYPL/L6ErlcEoRuhWCaaGvWL7uTd1/3k3I/
OMmsMwvUj//XcKStHoaraj+O74m3xWhyifgb+X8cEPrs8UpchMUcyi7GcXEEXMlMknLvheFBYQiX
OzNRj+P2Uog6whP7K9B3HfWDdc90dyadRc+wZnQFGhrNpsj1lW3HSCPivEfwyB+h9S4BwiVhpfeR
COaor/p9mJRfXR3hhOHf1ZQ3aD/guVSPo/mcGhWi6GBOIG3+ls3kfg9uld2sXaK6KGSpUdEqe6OW
h4FkwuuLq0Q0FkDL34hbO8JhO54rBdREiEdlerW+QjGt/ylA8rcRoK8XkS7m2mvk+iRoiaIWfKiB
8NdRLQwQWwmtuFM37vBzEjGMV+6AJ6wA8pKQE2dCQusi8Ic3UDDqsgi2JwwsFCnyPMaHZrtG6pGY
DZlATnRuJFRpFNRJ9JYCR1UeJOoXz4kcvRxkoTXHjCWQcHqagCmm8W2wlTdr0bNawzCsAR0L4MA1
q8W5aNCdkc1aJbi6TybZmLcfLficIyAGglXqZZPTGi+xngqFTCeV+mk8yG7rPnpI/zVwaL/sKVT+
37Iz1TlTBkLjD33DS0hqgYoxtbAbXwUhNOwr4qK4JTGSpGml6bMkIDpNfjQ/C5B70A29HgFK8jQr
uYhFipNI2JXXCz2sMONgjccBsRIWe8UdPXOWT6/Z+xS1Qs9FedyY+aejn2bmUvH0Fg8v1NLpJp0U
KMY2rNbJMuOll+LnUUYHuuu27CSMaVJ5NiiToj0+X12kYbBzCQK81vZAqmMFmS9daN0Pnbzqp9MG
XkNcuBJyhTGDfbEFY3bjIsMG5ElUsfWvQ+rhhFIJ4a7RNiXtCZOMZPcxYOb1lfJgmoIgKRe2P5BD
zPc8B3CftyydWr++ysr0XFcZ+STIzSV3E/gw2Q3rFIWC2aSCCRbhaBH4cdbQ/g7A7vq3EPtC51XJ
FnygzP27ieTIFqvl0b1gh1j2hz/omrmXwsDdfd3eJBFtkZAY0/ZyDYn0XEC9jQyg5y6rGWBd68Q2
l4N1sJTYOOSAsQkrqEfyeZ+XyaUZqm+8d8E17rSFO0tT4jfgAxezfgGdJmuQXkJllKaezLJza/ke
y+BA5ZVzoSCJSTK327uKfxqEes8cHgXV8b2rj2S5zYBIt5g1fPD+S8B740WFqhBQnF8qr1f39Qyq
WRUIzYA50oWxtYKSuvIUYJ7qoIIom3gs/lQg5MO1TwQtqKSU+CxENdz7EADnxxSTuC3ZUVW+SkBP
kp79x3qpmp6ExICMcp8y9LIv0KtGQl4m3vEAS6i/Ag0vP2n9KtMrJRInPhGpXQp80jYL4HVUmDkZ
uEinrEoX5qGzukL809zd0BxIb9Ym8SQeRlM1ZlqNdn5d2f0FXXv7RWSGghIUPTxMxA547lmEwPRV
IqkkeJmIBeswNXvN+E6Keay5WhSDahHCoRTKdjAeObF++FFLuaPzeWYU+KnngRBi1Lj282pBm4EX
A82/UO41pkjsHvHUQz9AxxpC/cD0M/UVNO8m0gUUW/ko3HhQSpp8w+iqsgVq/tGmPdRm5R6Jdt+M
PX/vCIE1rVewHYUsp7SfHcP8TPD/VIjrOwMmdmGNWdTecBgEz/VWUGRIiZTSl8GOxH2waj6NvxSf
1yp4awVhV1I7Oxuy0g/Nxou/Sx32xi+HPlwD20qRPjPIaIgxHByGdECL+mq9gazgiHWh2ixSEat4
WJuOmpPbBZvJaLmO7KUFEejsjkprvYYkfL//p482RO1r6YA1hRm9NiUkCkShwwp8EJffhdTJhs2O
xpOtk7AMYd4I6tkuKps3Ht+I+HTGklqYAzIpbEhyaoioNusAcH1M3ay+tVz/6RTCtaKSao8MoYo8
wEkEsvwYpf+gaPbcHqWOdclrAQ7J+ksSv78ek2exFfwDgKK8gMH1YhLCLwE5D2n1Gpn8C9ockETF
Y+SOhNqBZIXamnEEbjptTq6V+v25msS6T6C7TqSDbpgAy9OBuhVMDv87E0NhvladHrM+u/J3uU+o
MXC1GCTpEPu9UdDxf/JzFib+RZI9hb9ePvT4EwMNTk4632AZ6nAZQQqnS1TLN5Q2mk3ALfwIWc+W
ar/qWxMwm7aMsHjFbtVWIDb5ItNzUKQTNiRfTk8tSWIzo9FyO/wGXFMRnk7JCqb6bj63SAIzmatE
LHDglN8vrAtkFejNUXGEWzLtW7EgxNTWKhhwgfZGb+tH2hhBWC8ZAKlfDP0ym/q1EKc3UTCpIC2r
llmP0/B2M6jhgZ+n72bL10JlQHvMpGYI/Ox+TJgz27rnIrMehiiv/mpe3N6WaqbKzjeVBdr3If5F
+2wMsaMlQ2FCwzVrKlSqgcBFxXKGiOGGvGLCMh/W8ypXvXEBYSb834hcLr9v0DfJTAzAIsB6sEzN
HXstYk/xQjde9mz8PuhyFABhSfWDwY+h9XXWOCnzS4vhWldbo6DWpDSkgdUFXsQmiNBo3KwL+D1Z
8npv9RWG6PfhxkNa8NG51OLpg39m9IC2SeeLwSXFeFOmGqx/V80w/hexO/1hU4MhZlwK/yxaXpIh
35jrd/nOt32kYw2H6f3u0ImnICLxqwFDGZyE4gagYG8WFsoF+CxhjQHHAkFqnFq35S1KlVKD5Rv+
fX8Q7RJyWowPgdLcVZbggWq3y6cO3Cs85siKDPZEN+s0Any3bvFuj8U5U/hAqf5NAIcXQtkudPqC
FlCXeF6jzjxPZLRarEICUrFFSkeOwa6J2cuWubjFeS/ClQC/hTy8RnEh5P8VmBeaRIvUOUCVs/I9
EoVz4H+0vgIn6NEFmraVQW4RrDjopte3TM1k3WQIVfRcZUNX8Eqafx5ybPaf2Cy3eMcE/1MpU+l/
a9bxA0E563DOuqmmOGctfS7O6557z/MLdd0+iVC/6oubLKc0gDcbV983MjNrTSp9sXNyArGRYW25
inWzkpaNufDl4q6x96bQlEU3EH/L9J+Q1/yRqFLW8YaRSdEETH+IXMjoohWuCR3LBE7vd856B7vU
u67oKD5Hz7gsBTCjSi1cdMFX89XUaQhNRYj+qH4umDKTSdO471WYQGNCOnsTM3fQptxvGVLZ4HLA
4SfPL/OGz/+7ug0SiL5F7AWcgGaDuvZoBKZMeAF4B5ERiy8mAQfcE6YlHbQiN8lA9jMeyExR/nTW
xztsSXoPepNNEHv1B2heIYic+5+deL9pll8vL4fMP+KxZYzeR6U/ngntzdFF5FtpQSYo1dJSOi9I
HbCC0KGx+gTsXr7mnCO5Wj4wiAT0JPj+ZN4q5VUYHMrVIGoMpmOQBV8M9Zh9h6BpAUHj+0aztmFI
imd6x/hWa0tozlZ8pDmxFzBlGYyCBZ+NLeVcUcn+Fgn3gJuW8OcpZktvwRh/0xpaXtERijAofKV+
hDErracWCheG4eCf5fLZX10An/HkcQvL45Yyuqyf+Q2NQ2dzT4Def5yYYfNZkn4hIL9PLlXaA5rA
0lYqwN47ZVkqey+X+SDjy+xBzuSEdOD3Q46ZihxipyXrOabp2+OBVH6sXoYglIMNnL9yijrTrP9P
MNzHeCTAmY7hNPHt2tjiV8PVKauTpaOrIRg1jVlSd44yLWyzJjOReQgNAcsMur+Ld0ppCV62kyiS
jZP8ARuF4a2J23ojFTGsaUF2GnbXY79ZGRf/FwUVCzh66sp2u7SMsdPt0pzyfj4qTZ6i2K1Doko2
/QNBLC7LDvG2nUWMNsbZaKxmF3+XGZKI2zndTpRYg6bbR9vOSXSZMKEkHj7p0dZqSrAAcslr+H9a
UazxID4zBfXDkxEdxU+E2gZjHRkqEnjL6rKaOwrMGfCZurmxW2AJ20k0JRoUIfaeYou5XtP+cH3y
Qei2H8+26Cl1BI7xMWB2+zmzGrPDADifWNIVFsTGYlxZZeWc5a8sa3Ptj9NZO3ASew29gGXuHNHu
1H+5Of2uqg64BsxFXq/OGlUXnNL3d8LAKZnfcqVroF9j4nXCOfaOAm02v7jqhQqgo1S6ThwDgZnZ
VNyNHRmgG7YJl74AGvA62NAvYqyZ8jB5xvapNc+BdqbxjSu1DFcl/z6BJPW6uRfnDuCMyroqlZox
X8JKf0e0JYNSTr2JXo5zfEmBi96XOSccgy60HCzdm5oCdgV2/QZJfPPR/r6RQGiAST49XUQQ7v+1
0z08WxTYlBtR+k5m/KQZNHmViBVvj8i1joBzS+4/yHcAZJkov+DiWhvj12kwGKLGvrdeojPWCPCT
IPD4+FzSsO0fN/8+uoWypI13e7aSOuvoLt/ZjvUu939odbvptYv17dlBcU/vhtCbZ1AbqY6Tmzn/
WZN5tXfrsbQ3So7a9x8lFIvGjglMuebiPpg0dccBYaMzgfo6Fa9EKyWO9o69JWABnfxUs48Pdmeo
b0yd5R6ZcL3XSqleL6JcM2+c/Mwqgys1VR7Lsc5XCOg/K22seEiaiMWyBQ52dx2aRE63N3whhs/Q
LBtn0buSq0K38zXH9/076e0cErkkGeH7WvlAHDDoSVeXLuWErVNCj8H6//6Ul4vC0n1TR+iPpvGk
tANBikYEetjQDpfKqb/7wEYlfYPGmahPGQYWUBqnfEY6IxsyRB/Ii4j7pNKF+XI3i4lbpPW4v5MW
EiM0WbOZPjB6CYK9a5k0vRgcf46j5sBL301FgBvOz9ShB+UiVfHwoZUA7dxuMjZaqOl2h9v74xNC
e1B+rj6OX2xMM0kjzERgxsJKSdsK0ou5mKruEbnJZ2uT9ZdvHg7XaN+2W83WVi1CtvGKgIOH7Grp
1wj4AgyG8mShUrpmMhCHf3qRWFHA12VLJfrPYkEVES0ie8/NmSaJDg8jRrESzOs77rbrajNc5jdn
dnYcDfvPR8QdAzAKwEtPRErQeRz3Xnh2dlnhlZG/IIs4cvj1tOfx61W37JDXIwfpB/GQ0rciAnXS
z29wEaF+ddkF+LV58K0b8uDiX95Ixd42VOcrpVqfZNl45rG42EXHNDyHO8Soen4MA6MokPHAIaxG
S1FFnBz5MCY8x4ZPIrBsgzTeKbCMxzaD+aVag/Flo66TycJR9AEwYDiJSNULNhUBHhAQ/57aFFCI
cBLSJKW05hoqFg8PQOMQtGtKuOBx60VHZx8J/j4n5GM/mYWdPuji+k5RnCtUTy41y3HY8P5Sex06
cdcbr//HaOw2zlc+CyG1lKajXfe7G2/FP27wq4UZoxJBHl/ZrsaS5dIf/C9k4wVkeeYQgciU+Gzl
DQEDd4V+AArsFZBmVxs40CVVf0vACL02BLQViE+/AgBoC/89j2RGNzQi0d/JgBkPTeH2duVgBMXb
dp+QiPS71tW2wLBuREDd1S1MkAMJElWR70CL7zg3cUrofBPnTONZwlDenwTsPJgicbP3Nbe8+Y3r
oBONZlWr5zR6k0nIOgkcqifYHclq2H4lz1brGL6kWc9NH3PKayPv5JkjYhoHGt+utX/G4uZrNXbg
qyw0Mh5puqNubNEF8K5YcDKevG/3jwTsRP7yhJ5w0if5AVWPhSKeKl1iXJrJX5/QMfERazd8lWyK
ac1dexHhmTfO3Jar+Y2IyaWsenqsyMYg7CljiBOvNKwVTHVEvAPf8Gjv02DAUZQsAOjJH71SI6T0
eEUlm1GvMBKAU/VvMJlfMzjpQkaPKoUqg3lW6+Ah48ltMlPYa9DHteyYO27eJV+5QFGWhyjdBnam
hqie3RXG7mJ8CG0zgVg3USwVeiViyXbQrNbWb9lqykY/XYT5/SbqNLficob3FhRpFK0GmgA0I59A
jfVkegjZ9WDskDM3ddOaWUKsD12LwM8+IlYxWHRrN4eJNR2KWZXp3grOmqnig+9D9nXWNLPWFovV
lpIOQ2rG2mUeFtgPaDc39psRhxSPOzA4D9Mkm+wWhjTBYvXsg2S+BBEceKUHomZAOWOQqhy8b0t2
kBQd2Q3JzbeQlFrP6WP3PSqTz20+VXIp8LrML2WCxEyqphjoX5d5xXiaF3av0/F3JJE0mdFaKYL2
1fBHNvDMFqypS0FQLtbFMQkgxDoxGRXr8cChq0R43NlfpkGAygM06f+vkB5kCzH1vDaKTz3To4J+
hEi2XQdRKPaWp2GTgocx85RNI4Le8WvtfTxHABabWaHjbGCPXsCyyChcG4/VYp7lB6Dia3jomJ0h
iIRvS6heNGR8l2Wv1JyurdxgPQc+7EyRcxuZDhO68jH/WvQCI0sPVq+1h/8gQDqD2t++JhzWJ/36
+e090JOUQps8cUEW84+t37NyjexumIXpMjOXR/ArsLCGrK6DDbfJhviE7Jg+cnOKhWGXlmLw2WoD
2jhc/u6Q+hMHeN353qGfuJePb4bbaXdWthMgYotqdAkdJJmu+X8ZyZUUf7SoE/J9hc5kYdDfTdh1
qJ5R49kDx3R4UWLmkd9J1ZoKyg5yYG+YGJpqXf2eSgO4AvkJwJ6FBG/k4m1d3qeK/9Nsp8hKL8RI
vw2JFDsSTdJo8Hb0i2macVuQ+8ocrQylTwiocW8++J6N27ab18hcHlEiXpbmX1OHcSUyzo75ApSX
/eRcCF6Vs7C26xs+Y33HogzFT/eovC5fxkqIgeiSCTjHXZN/lw2T64g3zEm2D1JqjPpbQvM4NUfh
JWFTOiE9nYBi/WnYvRB7XlReTrnEGCc/fo3zC67ZZ9ZwG6lrrTvtHpIk+shgngyfmYCT3uxRWYXt
ybXQ4Cl736eKH6ZWKLd2aDinA9bWNbbwUgKkbUQlqzSM41X0D0g6a6IgcZtGVeRDel3sDd8jXFQA
qm6nqB7JbrhHdmpM03IJwa/jlivX6Dm9ghvku7rLjeC3F1yXvUK8ooCflgQEFbDzb9DKf36QZcho
GXzX2uULYK/O8Jh4EmQaqT+2e4r4ygczLT+3fKFBqwWibM+Fjmy7vPtIrr9WahSONEGvbrlayauY
8cG8KmcXBGnVX2FkjZJyW3eKdEggtMAHlb3+hJNO+qaibL/Q+kvb/E1caNWzs+bt3eaLKOrNNQ+i
URg1t25Y6Y2LIf2Gfx8jHUOll78rWUMl4Sjgg3wlE78gXDhfQPZfb9jOzpWZaRgXebCeGli/wGPU
1KqgStw6RJKmDq8HPkHmVeCqooji8BZJ6e3kJl8tNrUVtXq2nbpU3EknZgN1LN8KHtISfWOnHHwN
4yqiFd2jiJ2ho0urOsfkjGT846kFk0WrMD/ygUdVwFt+/vOqSVlE86sX/GNAsygJwl0INyE3GfYc
k2aS64DJkx6xAlBuNKYz94lepP/wGw60vgjy5v+As1Me6jdp6MV+RTOg2lSrCAi89Z7A7Njkqkfv
//8qME/mmGcSuSrXhnDifXxZs/8eZT6l9qcI2np2SdOPw8Z7bztUNadnR0fLMDOqR93kKlMGONPJ
p3iFSKgY9EbBBsGETPrMAiTF1llwnGScXZZdo1fjJzB/SliwtRYMVK20tdGA3BIQ4IlY0LDLY7n9
eHN+/PxHLl3Qb4amzkvnafkx8KdkS8FzrGC1zG7thPOMwDqWSVNl5rVSbkwpZFAauAIeOgiFivZV
wWH+K2rb0IVmEpgkezUT0S1LgV5S2d/WRB3BKn6dR8C3jgnD8pPqlctyB0PzUXwBWMFJVAxfs3dM
FcE9R7zMwAwksyFrwW81fWJfIENjB5DDse2m7ro5VlwzGer4bO8yFUQJ5SBG1F5pdgDDPMX09ci1
502c8de3KfcevjST7lFUTvbsvcVwVmJpDCKcabKjwvMbUYO3Ky0uKPJJGL3et7MsRkO3KTNY0XHo
dNS0zixv9VQ/tSdKci2VPpdCel1DKiwxtJbxeJWDf2cWJLyHxQiq5cyXhauH/qyPhvvPHFLvK267
h7whYK0MudSH5XlFzpATLfYRwltVF++yWezOi0+vXOC5JkhmYn75b0HarOYYHiIvCokwXjvj404l
VOA7cC5WnVeF7dIUpAPeV3vKSoG6nwGtG5ShoZv3Vy2MNyngleT2c14WS18Cps/zUBgzvIvLzGra
NJTt+6T9HiXRIxGn1UUfK37ytOwZ6IcCZIJUSIOheHZuRKRqtuJu9VrWoJ/yxvAPPLLCeeG3qbV4
YF0KteuCWqqicYdXFP2iHouWicCFWJ0L/M3/emS4fzYsQxkX4M/rTdmmjK2t07z4iHxNnNvwpbLj
P7ggjiq/E9ZGnjBvnEcXcwHl7q5ybyfw+906Aj6bZ1SmAFYcPD9RvFJ5Mo9f6R3fplGLSrKJiLHy
St8YN3ss874QHYZ932inPQrQfXPwSIRo/RcApOMgNMHBhB5LqFaO0oqgrsMt1zfvRDyOJKmqeVk3
EKn33tg63cOmv0d+2a2BvVAkBurCYy61HYi2zlgDf37jM3QNNWuf7w4sWbZNI1n4rDRGJyECF5ON
cK8euuFIoSClyzi/1xS1RNX0msmTzGcStA7b2qifZhCACU0/q8+shCncDculdbNStM6ywHpNpVV0
auiag9Rj5DbBXioqEqdpTIS1muNTQXtoYOP6mUoewcQDmIhUNwBo7KwCE5G7RL/S7NM2/KOEVe06
i7feWVgbvzwWwNpVvRM2o+KbCqlpDPn4Hd+hVfs7Ct14t3gLvxY0i7X5xG1tQWFhEeZl0qG/vrD8
6zIOEGbdTl1D+kHF2uyleeF0cCf5gxhgnx6X2N+yiyxysyHgaXAF4N1cFMJ8b/KwBv1sBpteqwun
NDjyjnZdII/Icx1P0hyUYjYg886Dui7+VnxPkBKJX4T2Ng0QpZd5mtITMlRbpntFmw4y7vTtz0m9
oj0c7cvDZKYlltKec6hbTnmKYcZlKhLjmmoAv2GGMpLlGljTKXPkcCN2kc5IY7xLQODQEb+O9S1E
cXvk581xHzq7OUWeDACTl3Eriv6F+urXNEDnA3V3m4fKjt4UW88MbY1FSeLEF8+Xk07V/QZJClgs
SvpisvLpEbcNNZ2rcQnU1n/S31s/ZeX4FJqCe2dbNLTrbqdXDcTlXVJMw/LVmgcoxJqEne5xp0ig
UDBX7S415A7apeYq45SmCDXlG3JzIcW5clvwH66gZ4MQjug97idEunwoGmW8FlyJVKHO5JP4DTs4
w/4NgSGbuYM1ucHgpEopuBKUlkgbEFra1Svuyx5AriTxaXClud7dZoAyrLW8ycirhnXFyGq3j93F
jmashzcAQ1xry+cAQThGv4OgL0D4ePKwWSHPX4h/0r8/uvxGSOfAfgjAdbxWBRdzqkGVY81axapH
f+SKBbnMZ1GIJdwpaNsHDnC32lAciRHI8PyEItvJpV1sFBVw8Y8d5f+ix5tIAclilgK2oBz6yxdS
LnadXJXr1OB6vgGWavS1XbLUttp3OffmrYu828zUmsBFDXGXVFj9woSaqBSK9hg5YuXIpCEmOheK
jVdRqNBmO+PVtBIfAWqtTiB12IT+KW45p/yk2INoGaIvAsJ53jihjMi12a3Yux+OCb1xPgsAkSyU
Mde3rNR2VNW1Wfes3oRhdSW6Mtvi5hFr61cB3k0LFD/L98rfX9ktL+LzUOd06FYMJZGFxG+QWTbC
oclNpfT8+O80Sfc9b1aEJtV4tz97IEFvQA1A3ntxsmhIEgQCsnEFCFGtsU056KAOQDl4y7mbskX8
5DiquCRgxk/QWaUvX1VXuDvjKILrWpTix3PpeuM32RST7ljsE9eAnlEf5DOlP2f2yUF6ik9CsPyM
XLvp15U2Cxoy2vXVJ9wwbKonPHEXJXRAwhui3WYLa2chqiRfbmYqMe214hjDxu1AkY4wfeb1VrQD
NLPToDiJ1o2VuQ79JoTTPYcodcdZ5ug0yM4QFKiii/Yw6GqEjQj1HyGWzAOB0sVb8GPItWFjl0lM
9MfZmYwmqhVpNBLskfYReEUrjHRdH+CkmQbDeZ3Tl8ZXvtdP65CpyTMb59v0FADBhfVk+aAJZ/aM
StiWKu3Zwl7i3IRWA/OcVVGSXm/sP6gTDspTHPCKtIkffxmoX3UMOaG0xuj5u0qIXOf953Ouwm1/
JemoWGLyrRmF/kr8ylcpgKEj2jpdsYDS6XwsI9CQweZqNHMZdgBoMyXZO4opPjLBb6U8skvNXOS5
OvrwqmLS9jA3S/Jth2hLLD6JQ1lmCoNglSZwx86Tz9zAYqf4DBOQMdbK2qSsr5PSWnNtyKRaqazn
MJleSM/exfKnavX416rMRsLUcvos7u193nW/tfcTdB+BWbcFS9XCl3xczAqbuEFhspHasXFduyfa
3F0HUfutZrpZdLWKdHTgEeA7xqohoKKshk67zvlth1jgRazLOjwzmV29ADm4fBIIPRgV8Dxow2Yq
sqXCixhc+ibelzYFc2SpFLavNcTBe+wVFgbfslPiEknRHjTzGqOipY0a+0YWH01e1ZQZN6jO0oIZ
kj0+Rx1tOZZMVD1UuMNWZJ5HP33C4wY9G+H63IGj+PBC0JxVx10MN5ZQx/c6p0l4RBXOpwY+bKO3
dFlhVUGrfunBy4QYEY9Zn3FTC+RlSmuw40KPhLbkcERjy9nUgSdC+JL7ongmmzKYRoaiHxtLAavk
KktHhYmPRAYYAiESQB5T6EyGurqx5+PFjQPmwWbHrA4x74Yz43CcuNoTWVyGHJ1gl6aP7kj3wfBY
xSVJGs1DX/o3IurqoGK3weyzHChS1KHnDLEJHPwxESuSrKPGs/iAurhFjCa0b/WtLLwlMH0/xCeH
PQ0Xi4vHNP+IWJRNG0tAYYo4FGtdgKNDxbidV65Lnw8/EJ8YtrlqkG7G3yqC3HcGJpWJXAZNyylJ
FcJqGHZYnm+oMk+jkn6mdHeFBYJx1Rp7gw2D4tmY3wEBrmRI9bRFRyoleqTvAhCDbaDcCHlPlWxc
ChqojpLfCvIHyTznBaRQftXtnI3IXq2ET+RO89Bdr3l5V4PRfpCEQWWJzQgpJcxuctT2tuG91XFL
dciNKZ3Fk/tI0VfHoxgKDGQxuYUJEL8PSAn2qsz4quHDU2K6xtSKKkLNnKquUWfOELoEy8orjo61
5RvkyP3LHNPvcaaurBZSIZ6OP/UZUD79gNQPDsi689zQwZnPqzlX8m/tdzmcg7InrEEwbJle84U8
hlK+sxAmHtN0zP7kjLfQKJU23DcpGoX5Thnx94KfqQWp4bZlWZFxkHjJgkRKloJljLZGMoAAnrkV
jrPqrZuv9EPVg3vpiY2Aax7kyKBtepW6thSg9u37Tj3mdR7GouuSVFjBco1G2tz+W5UDki/9yQ3i
HjdwDXzJm3X6rZiuQs740ocqvfptMbXWRqS34zfv6KibM6S7RwINIyAJUwVI07OE6710kykb5C3h
B+AKEPjjWGtpMdTrhHeQONDdHEGCd7E85+Kfrcmwa9X9Te2m92szropkODo7mLy2BgTrJ16LU8q/
C5p3wUHNU2iB1/Xog1e1nDWiDiH8sWViQ1QL0IcFxDH+xDPtZUVlCGuSorYCpmyZuPfNePdk3qsd
tL/ChI9pOsLGOhiT00DkCM4kKgs153wmM+Q6toDDMqRDqgy7oEf/9Oy14teArw2SG0REiHDnktHV
bISSL4otlHvnyojIKBvSGPKsFJrnPuApwfuXam02GxOOZeGmU210o+fJEGYz+Cfhccc6+992jINo
UURb8racFMXe4cDXOx4E63JPgD40owBeT64CUX+YVQj/5tiG3aWYvUsgGgwXw489USRHezjjBW/f
cRkAoRfuUoaheSJ+qYYskhd0nCxohRq+Tvl1iQmQU1xosJArZkDkJcj3folkrO1DDxac0ia8a4ED
z1z6p7noPJ73dwBXFmvsxq/mVQctcah/IEF5ERL2Ymt/yqP/Fu9e/8Uk17Ne1PrOP3ifttgkJmvG
CXpAJDFcAc7aRCuLs4QOqEl1WJK6UCEktdz3+Q+i1TQnffR6JWVUju1uBgpeK2V09Rvd8X953KiS
8BhSzbTV5OaaZsz1rqPgEJ6axARE4P23GR17G6H2ZHf7ACUm7JAx2f7bx4oH89yctPTov3iNWk7f
aR3uRUvyPq4GIKWX2I6OxJES4dHE/9BnY+wQMHSfZ1bo7W5VV1sJb3S2GDjWr08cAhJML6enVGJ9
KGhiBfQQruKo4Aco1qq9U5wcfAlcyfpmYk4p3Jo0x8pnp0r5NpToYog0uqa+Y+wuIEOfdU5PqdSr
oXuZu6M+sT89ADufLth5RipAcOP7GkTGOVwWCUoMZRF1i6CcHH9wNGx87WGkqawxNeEPdD4X+4hf
wu8BX0fKfB0IkpP1v9Q8Irir25Adth8RDXeWMg+vvUCDb3KidS+pRwFrexTFhFbcr1HXrM53PBUG
psOeZlu510/YR08T9PlshyWntEEfNl73V22aznZkb9KfWObmaRSyKFN42EmZ3IhYInhX0iF5ox3x
1IKvySIprIpbAiv7J4A6NbDh3oH3841Qfs8o+d8bUoS4o61riEeFBABzKf5xT7pXHZW/sUu8aEmv
0duhGIsC7hHaa6HolYV5rh4vrW89WKlaVk/z1qnw6LKq9xcd0Y5x7FI/7D2/p5E6d47qTIDTUErX
CaWrWf9fT9db+UqaNCwzGFMz9hA5zJyyvlbICuHFuqWV9j0DQfrYj+4pkNZSUNgUAHdMSL81cmVy
jXE3uMkHZfIzhwYgnBz8FNPNl4teSg9NayF0e6gZtDN8aXnrKHCXUbB/ubpef+vPf9g7sXOueqyR
GuAXsTtsXfmNxdPtaXVSbaFSt2YETX9RwRmMjvJYaNH2UH/2Wik3JBma4cCs0PGFIgZuXH0ycRkJ
iswezhVRrfzfWmM+NwJLr4HpyGqYWZrmIiA/bTuSd8hXEjQ+WESSbj98bQZD+iSuNOl5rEjW/477
RdPlajRh8jzIrbznndv67nna+o4INWvDiyktVTkTuBpT0hdDLxegfSF5SHPH8FrEfiULI8h5SjuR
tFs0QS68S/+keJM82x568Od+gReJXAa6bJMKVZX7su6puFW5+3DxGWJyxrBWe+4df9fZrHkS+E7x
e9d9xWC8t7DLp+16gkDVP6yGSo+lK951KPl3nHw7+aUEF2YM0PgPFPva9/Pc+2i6277sLYaPkdIG
d3a0GYy9qOLeflK0to4AqlyCRKCc7cSpR6acH12inlD4tUaBzENGQd85ncORBQKXVJ4NQNzSrYFk
7kM4yJicsCxx9Tv37vYW2YYgZGzgf+Ta37XiSF/MxMg73yjKSK9qMlg4sdS9sXNoWtahEtXyWnlS
ru78XdlzXukuFs8tFZnjHIRwsRkuf5CcbDnKkjwl+XvMpWW28PTy8Z6gml96fIycwWWmXqwdX+aG
Aw0FHWB28M2Pne57rG8fZlqkdTGeRKskSLtAnAdkWbnFsIxlsIq+mDENJURrHgkBNXAd/QDa4sP3
we6LE59XCawRp5U/Gzgo2pZNWAeI24FbMSVX6arLyIHuw1E+gNrC/HqlmWTnF/iGqAz/0wej9TQg
IhAan4Y4XGeEDa95bfmLC7eDQA1sna08hyhm3tm9RdsIgRTSRGMaOgIEwjd9nVC4CZTP1MqI8FF/
0npAA9BRCbL1hchLG1HE+JqrEyI2czGa7GrcyDQZ61GpA3gS2Ysm8JjToAENMtDWnZ4dgYM8tcHO
sXFyzMcjfAb3cd4kM5O4CJcGfD77Xb1bH4rff+ft7N32Mv8v6m2diufNEOle1HFvtkjqt9nt7JcW
dT4mHCznGjo3ZHqdQJmIQ0eiKLbpGTUSqaOAgqXQpldJ4u11lwSuxYKN0AuqmmT61dzF4KMjwF+b
8kQkim426oa3snm8tpwb0k6Nk8bQBMtCyRcZnr81EMNNUcLl6nAp2d1oo0zLzZqw+owT5KuThPhx
51iHgx5N02KnT9pYiF4peo4BFrTfhRpQOXofFaorMg4su5I22/TXomkFMxt59mvkzN1jbRMfYRc5
yuwu/h+V8hwacNSMrp18GM9ww1k8CezZS7x21jEIhuhrPmwG7iGjUEdFcBtdYoYt/XEx0ohoSMWU
Yte853QfiUA7hSgUTE2DhLGQEXJ9lOj/mgTkD+3xdNt1I6RDn2eanJ43EQ67yceIpoincVtXkhjZ
Yxdnxx4+lF8cFfO9JSzV2DxoAXogq/iUGUrDoFegwMs0cuW7tNPs2bsJQ72i7Gf1c6tqZqCIpwIF
jir2LXeRbkXd4eSubJdNEdKHhJqYfFjlQ18BRQ85wXy8FwpS6JiPTK/zQoYlTfKLTLHWJ5VqcC1R
dRxnRJrH7LhVFavK0/oF2qBOzltZi4OolL2XYLHcFzD2XlYN4+MZUwfoc9B4wIit1dRa+YPnrdKe
KJQZ77SiZj/hGRFWFIQDYd+409eC4BH4d7tebeYKDmdVdfTj2czXvVe1pj1iW/vQISyXIk/Y05QS
VAJy26eQa4jFam1BxJ9pENfxk6PVgexLYsjBcb/0NQ3lMgtC/ktLArxD8RUEMp94WOK5kg+zmka5
2VTWWuS0HeWZtb+EkncIzheATOqRNmPAdpENgO+eBG41IOUc0x7GNZgBKYA+HPpWHcZHfiXCrdUU
YQcls/xmj2p87JWvJhfVWPP54wtNjxO/mX9Ig1/Zk9ItkxtpQ7t53pxInfPEtMeG4a+UyzwEpfIp
XcSJw74ItHit3Fd5fAXdJWhslYiPIcrsVWy0rG8GcSJvwCZGMesIBWgclmQaD0z5/37mxpBo0Fnd
2aLPRVcACnALvTTGpxGj/GCJglMZ5cEJ02suCzJbFWUDRYWy6IDF1h+gjrA7+lSvO91jnZ/9Am2k
fW0iMiABxO4+U5mdiVLUCLzXz/RZp1AGTYmV/oW5i8EzSyGv0FrUSPInvH3YrEJb6Wa9BBmI5Bhn
X1qlbUKiEz0+BNUmUc2tNg4hmNsVAo8XXvZNclSCVJBSI//Nkex7DTQM2+TEqwc/o9ERI6bUtYSK
HnJIJzvEb01fE8GOY4NPtKLW75vqQ5SmIeKCG6F5rvYHxQjNs4Az1/Oogf3lo5m9kjkEnZ9H4VeU
LIimilgUFsqfqKWhbty/0K8NZcGMOnQReaBgRU2rj8JzrrCCZqdXJ7KxPRjJZ65+nixMhZNtFfly
44Nj0lwQUWqBmjFHoKyFii/p6BcJs+zCcA2G5Ks54jQ1KI/ELoH2GYqnQBpXeKSQro/SCT1sv/4b
CKEdXIk842j2zdE/tBEMlVRab1JYQxNvK7EYCuf2jZBUrABFrbgCs8zv496YAPTo5ODUjgpXNv7A
NZNT7u8wmAofMszpT7XUlLmpda72iQmyYpujzxqy6o++UxjyYUasP5EKAXN8+b807Lyb9v5BlKhG
2fXdki3pL6oiUJODoOL4s6xIOtt7DCxb2cc30IJWnn7jVx0oUZNBd5ybK1g+fBHbfH2d4E1BL6Gq
NoaMlmcdq33qL5GCSG340wHm1rTIqR91+EVVpSCme7V/CPS5LOUYIDcEYdIRcEMY/gJaVyHkRJdq
ADzRrRwkIpgarR5Y8PEtWS8DmIp0LQQgqSYQXzBA8q7zJS4Oc48d++VpqoqfrFYQxbhMqgBboy3l
gNlWMDb93K3jpr6j4N41Jn0QLI91XM2EsX/iRcUpGXSJd65XJA/FoeVtHqvZ9KntX8cP74oB4fTz
YO3H2V26QOUcZcOuuUl8co71hPb1/uo/vWg5hD7OGyeLnSXry8NXp7/VkptGwR57wMJYHXbvbYhh
V7dMnqjHRjLl+zQRRnHVu0s7gxATulst3EiMNMWM/bkFdbYIpJAjT5wuAHOMwEhYOWE8XTcXa6rX
aFI62vyPp2BJRlr4ak0GB22rJJPcEbiJe1oVJpHuD2kCy5lUJriOeEfqfCgcjVddovTBB850/5nd
QYkohuhZ620SUjIK7W5tgDTpfKy9ldbrCG4oCku7W6SyIBMhGt1oEIFHMu8F0mLAlCHQzyUV3Ejr
eVn7xQrt09ZasNvJ+C6OhEo6l9rK1eHsy0y6kC+E1llvQ45axG9OLaCpU1n4gXoUG7le7XWO1Z7p
kH8LPOwTaLZL3hsSUYFoYZZV4iVmirCjYfsaQ7F6It/EqwNIni0bd1furFzo/78qWE3FYbnlFl1v
KZCHHnsn6YxLZXmm+nVmjI8HEOl3tJZOJPegY5lNEbySaPNZ4SD4qx9uo8kldH7Kx1as7fmGcDOr
Y8WgLJzI5MyMqOcnfTGeATVnV6qPMSbSJyg4zWYEhWQa+DdvJW/UiKGmWv+WEtmNOk71gmTL3gJP
OPOfi9ZqFOh+/2MT+UcFy0KZOvrB5pbq+Kh3ApdLoyPoKvGB4HS6G2JtgMVDOOWe+8FhdC0dCayU
SiY313gPRTVD4I8sKD+t1OPv8jGFWE3jUijC8bCOOHXi7C6UjqrMno0Lc0N/aQ8+39FvqtWJU6dR
oTVVCayPyvbKgkmZHvGiEByw5qAl6KxOE76hcDxrwYQz0sNSoa5U9aj2sd8rCGbNH0g2D4H4ZJEb
rk4Y4YIdWMUNvZrBxoJ74qfHuL6BipAfNwOHvUO/HsId7uxbYKQkH4lzaWgAsiVrAT3Nqg6SrMKz
hx3KqMLZ4rwTcQLHaeg5WNTUYtzzxGqvzqggjDrEznBP3bOm4duTxjW3oFSVVyFAQbdUuXUyCWAV
a9x8Zqb0Ac6ftuRQJd2sAYb6bQ1458vWwJoZ3P1QIxiNlMmJKbxUNJXksnZRY5pPK3vAoOPp3tvC
oZ/dvYxlgsXjCO10PBfLZdkn2yjdh+gXoOru2GuazVVk/zNZcuthKmWx0OIUCzMzpuCV4DTm+AbD
zlWw6Z0f7+cURc1n3BWM96bX+2Am2EaKaZnZ7+ggOYlz/bFAbh+9rWt5vV3aIU/V7IWKcTcllxMG
EI8HUa1KM5yyA/QEQ7YhlilqzMWj9qLEbK5OdBKyOMq3t085AQw2sBnSF/mZ/JiXFC+FZaa5SCEP
7Wghzof2IZ14x/dmD/tK0ezO3v4x+JGGnEQ0lVnGEWA0n9pcmEDpcBrSjtCrLbRO9HV7mhhm3mLu
8hoBtB6GPUsHFlNywpRso21G6D0sen5tewSuk1sR5VxP3Z7PvNk3GbmRxeApqQoCcEUAE7OKasCq
ckm3MsihE94lhpKuOBb4bLvQuePtqE5L3OFXXqSxDbXfAgdIcQBvkBMjhEuH0B953Vo1Y0tMaGnn
N47GhScVx0LjxWD0OxrwYgc9PLJ1OKbv8f0kprcK4+IMnX3nTjSue7cwEBcn7nkNVcz4SS5kSSvJ
GlUHH+YmupaQAWjDMjUSLLg+f7ZNxAd/GcbyWh2R+bEMuNye8roRb7AN20V86zGwtFE8S9hldzaQ
3HaGUsbCZejnMlagPJdN+4ydnB1A2bf9TSTo7eA5nKvALxRICaDcc0iUgM/dTLDPWhLMx0P37ODn
ItCwb558r0I7b/Rg5ZB1of7jBhdp9/z7daoxloR1zaxf6mcOJB6FZ9GNgiQDRe9WnQK4m1U99Mw5
iQXIRS0uc4esLIjzSiu3aG0mknXMtOtJWv34jmwkbcCDwqkk+vJyOj5nCa5lur5ATlsJkEGShIF2
dzkgwv4M3vxXTqmgxmVfovVkyE8K88m8Ra1z59t8MCZhTcvrB56+CudfXBi4lIAissGAw/qpfRVK
D/7Ol++S/0BPHOveqMkoys+dfh4Is9pHiXT6znbzlXTD0fJ0fqYUt49HteHuXhufd68EdLaSvzzn
/osesWMJDm89JCc8XJSRSmcftFhGUjjD50N/SxTloVKU6eL5hFqA9JJF2Mz0iz3K+5mGgEQsDvbe
tCa3QlwL+9De0zu4QgupW4qI4qpNbvsfGuLNBeJIFypiCKkbhJ7lpp6mpzJbwSrMXnARRdMobgWW
H1dlB/7NsWQVm6Am1jlJb23To5OTwQzMG2QVC+eQhqBPavUY5XXcy+TWysMKRmTUmaSPB/CdyACP
Brc5xKRCO1Q2za5ERvXy5Cr4fxxkqEwiChfIq2339J/sjBZp+0/F9xm1+vxpeoNzaGOKmEdhCOZ2
EyrJTQcZXhWvvjAuETBsilZ/rDlDuiyrQ9j7KK0iGqG7k42ALPQRtKd+WyUWFumuKpY1THC7wyMC
mtKj8g9eqbITXxPXwIfJzq8Tssqhqh5exKT+7c6IcxsJcfEslwfSep14bJPIHHJQl2OFaPSDATTi
2xjPsItRmB88mSnEnlJGgYsNEcHXaRbl+dxM7vYXrE/w5xaDQdMWBAm6gF+SYD2sDpW1OCxUU6pP
VRoSEUpUu0g0WUZdJFaJHeeaJGX6dXD3pCi+zvsOHFl6LQEqn8JrG+h0gTMQYGs6z/s5eLBUWZs9
iqvxLgFo1VO2m0fn7+pEKcbMnpDR90i5FoOllV5wOMGStV/Pqooi+4budubKGLlWxKUEy5LKAEXT
T1Mvjf9R5m1QadbApJD2MOO+tJuA77K0npIlvHBDn8oXHQV+N2a99BucC0MK+he6E2x+gZdxdrPX
q4BrP8Dt51zC5+MHgxuiro2nIKHF3uQq50vfmwaNMK6ovNailQXu/zSgMGN28FLmVpdIx0VRIOTk
Zq01nFwOlTDiy9qxDOQW1bSmm3xrCt11WTi8760D2J8aTxTX5syetJ2LULem5GzJT4N3AsIp25yb
YCKs9NgFeIxl0/RKO5jpag0IIUEKOIK80Hr3Tt5igei5vAGn64L4pbW8Qkfmczz1fbZtv2+g9p2H
hGPQqrUvM9eU7otJqdKXK/VPa2QTs1ZpR/0Na/r8nGoE13KQCzKhOqzNXe0kiXaJjRl+ZsyzJi+A
UT5Bhi4DZ99qu++OnjVO3vMqkxCKdswhA5M7yqnA102QlkFKVbBIry0I8LLrHECa2lYOaAKMHzhw
niJyiOSAEBL1+tRvVPlxCuitRQ2xZo52yIh/073hBiDc/JzzPzffzj+8+n8diYSaMFfZ1quRVkdL
QxeUPmx7JnAqTrA6UttJNQ2NToOBQFc41NtwQ7G+UEsKbQx8WDSq3pVNkWi85sLeHiUqxmq7nMBr
8IA0+HYLb21E0oQs+RhdF2S9UrWJRlng+fqSu22J9UKgvzLHjq73S/q58tfLt8RJFaubVrZnwwJ7
iloR2o+Sq9/b3jO+PcCjOsdRYeO7iEQCyRufpH9jYHzu+6GeCQMy7hooX96p/Bz68Lb5NS6WmXxY
yFktj10HN6ByyjHbD2Cwy5XKOkB2vl4P4qtE/Uz3vjtb2S3Wx/4KYMM1fRV/lBjclFK0ThKi7vb8
SuokOj/Oda9piZEcmM0GlnVpW31i+8P9Xw1AhEkWri10dr+bjgdpxgJWQ9FA3ZWUK3EmK5BqTx//
vRs6MheNGJwhJLem8tTJHS7OmO2oTVtPo+KTyWm6zYDvQ3ODpvHrcJD37danXZIbIhosFgakh6hG
K05l4kDnF9U9hxljSW5fUIfqMmxlwclJeami/0dKhhucNOA8OreoIz/erfa3tW74ouh4a4Vt4A7C
E2TOVP3MmySO3S3OJeOEmu40EOC3Knui7tDmlVLiJoBsaOxy4kyItaoPIrtgwWHRp0ehJHxf4swH
s1PJpzDTOSbv7lbyGx5fU5m2xHEPfi20YfAxO48AGyAnuZoXvdlKXHZnlsja4Z82WFfL2SShualg
W/yb1VFLYVkHyoIx8bTSWlccoLnMoarCP6X4KxstPV00eA75qR8Eqj3DOz0c70Y8ZDLo4DleAApv
i8u1Cqrv8+ASIcV8V6SAr5WLYUZLkq/MPFy+xLjPphktzIy5Ar7pUkhqFhqRQyr+ldqDTrlm8C1M
E3x9th7mfJ7pIDYLMACSqo/FJ4FxiJmFimaRracxtMN5Una/96ACvadelwUEy7b3QWxEsrDYYYrN
zRJ5UrQhkurnfYNDvLoGppyPhWplkwJkUuWTUPEx0c4YHB/0mcJCkF6qP0IVrSA++SQXbRMF+0ON
6bWO2sTaWZZssjlroLULwzeypjDGXV6yYEMelu2WR0fBkTyeZtR5UCv9gpRFmz+AHz6/nLaUPXmV
D2nEjtujf93key23g7cIiOBpM4CqabvpzFUMq2Hb4umnLDve3gQwAucp+5GnoH3dE1GV8/bDoGcW
wQYWt3EDp0ftuAvgSnGwmSNffj2RXOLPFPzobFfBNPJe5em1ut17YnCYQcT1Q06C0eoHSZDnbSp/
YIsiPNluJvgaOolchCuZmuCMhFVtJFHkzONBpKJJT6VGCyhLNyhmN1X85wdDlJ762GCEcynTWE+h
GqG121DUK+ZOEyXzWzhwBUSByFUTfdmbDuo89FjU4N4FmjVc2exDhxzx4AjaN3+D2Bmn4cEaY6Kd
JdLHDnzIkeNdEKtQ7R/31gspwxVQc52D/D0nIEkNfoKX7UszdiGwB56gl5Y6t92ZF/BEjWVqXj0R
uOLyCeGpZTq1UdiLRrIs+danWPJrl/HtYbhZdkHNzAwqgXFRGFUt6YWkrTtKkunB2V41lGM4IXXj
qHMtFNxKAU3+zQJ9Wtcm4/xW06VchJEu2OPzWhhRJaWfi5mTpneJNAP4tmeylWvAH3BfmqdrF1j7
3tgQvZvK7xjUxljyrapLZbO9FQiHQQUpfHN1Y3uuLwxMnNL7ybNfdP8vQ1NmVPUcJg+1IYu3CV6F
EGTzc3gkQLAiirw3uTmSAAjfsRF3cWiD6tgFYysHavbxze7bIkNk48giWECsRAQRdezbN0vh5mRM
Xan1AMrZB4r0bXftXHYvyU7V7JcBU4l8Mn0g+5+ULLPL8+nVK3kf86J2Z7EEYL6mjN3XMlA55JGg
russ9rlh01rofkR949qEf/QdeVIVIrXQOBiatEPZlRofWXg+SNChgrf2HyF/eH6oytQHks3480Gr
bLPTN9WsL8nEDpvyZJywHlfJUuJCrNs5lFscgUjJDamAP7GTtyCLdQZ2lcg7UdnGkCDKLNPQVwVZ
gaDm1ubL2lLGZ9uLbZ5k7C0nzw3FgtJj+SDJgD0rdj7amG1YQp52SPdvOfMSxtsUhtKv2fEOMZ1T
AleWTq4mYce2FpZyc1Ow1g+HTwAf9hyzq0z69WB+U69JQcd0MkH5jtahs2W/n5Kn+1WEx1uPWp7z
PblmyddFUNmBdEecih9tquYGktP9RI4I4RiTP57QeVKR3pzyrph8p4KzZfDgXWsMC87XGPngbTkN
lCUWXgzOOpPHj+eLSmuY5Zt1WZk+PcNPJHjFsJEYICXePX2xUtzjzt3MQiwfSXIg6jSMvGMqDZ8h
U3gLhJEwL+p37IF6cY8WyNQa9sOafU4SfbQP/yrvNLiuklH6rNvoL74CoNmhzVCU2BJ0gBJZLd+s
QXXH9QDctGFGD5kGOFHw4lBjmvBfu7u9P8CGUrOFyqHyJTQuAKQZGokvZIA4nkqB3zeT1TvwHdFd
Ur0UCU9rC9QOdNKeszA6GGKpU+ybcrdeLSPcSvi2k1outaN+I7misvrhTE7jlSagsWWDbI5Hil2s
/ILKQYNGxYDED0Ob7LnRSHj39JexFdVsNPkVPcQa9rLwDSh19LBM4m/s4hht0IsNk1h8ngYf0nsh
WI6mv0ovlPZuEcyE6ckbsZ6WViA+iMyaFju2ghLKTVUwB72OqCzWwi/LYSs3WwY+gA/079YrkMxz
8/AJ1kO5pohdP5SpEdPaC6B4x5Oomu04tyKWgi9C+Op+AYAyEf0EJZR02AfoQkHo/8dBudhxL7HU
eHUl4vFjiBBB0UpWIOhlbXZq4Lt6axXSfhzEP5LVnhBKaoUSUn0rsK253q1xD9/8zQ6hsuiB56Ei
Fprery4tgIq3/Bk/nBpsbNZg0nNtKQbq5/Y9vRFZwJgxeFUYh0qzg7DYFMNGARHdgYIBP8lqRumv
rYC4h7vJDoBNatZwaTULpwOycOBeSc8RT7xGp9+xXcFF8hTswHAe1cmzf5VobZGetMjoDOkz4Aut
x/EA9EFAV/L9SlW3iNr5pNtYIZiDVYVSTTBRPv8G6DAc5iwWf1iwmkw2ULECYtnKTltJcNGSUuak
rJesBpaYz3nyy1GtiNjJt169FGc1X16M0KmxqaYvit8xLcctEkTyjf73WsQT+fZUd5V2oMXm2gP4
ykMXKqmofyoGgDtH3NEnBKCof8hs9OGmez+EJIhBBhiPd/crc77ccHuir4iI65Ip7MHzvEXzmh2/
Hkxz2ZRGfsnZGl/sX98QL1/1+CsS9AKzg4L0FJ7h9uUqaQL+CxJJ0KseobDsLTtvD3wfnsnocUji
d9p17407VNbYGIGSqls8Poi2xwetw4+ZhUp5/oDTqbofldgnLz0pI0vZ8QqcB08cK0yeu6lGHK7s
miFsntyZFSs4/RobMlH9mHsdEUcA/DdHuCT8Y+Su1BjPrTKVwxJQjl6KrNW/geF6xG2RszGU6c1V
AZNHlLuckV0RnJc1Z5ADC6MdCkWjh3aLAexsXe7OoSLGsMxADXzCiFAm0xntE2H5pghOKIlRUFmc
BcWy66DGd5FCIAW2kIb/qt8VBlJDLhlu6t9yTI55zA6f0PgPIjq0XPnRoVEGjLR+lrbwyHaJkUDp
I2fow19KGBsvBUe9YYcyuP2MbYHosE8SePtcZm7ffA5IwqOixDGBKF0Mf468Acd//AZQGagFJH1E
97OC+LKPrTurQi+nZa7yqgBeQw/nPblHOTYV2fkww2nIKBMkhxyaZg4v+9FIjLfdqOZ7DWj/GJV8
jn4ULomv6T98Dw9clg6am1yO1vKhoTBCst4dReUSR/CUaYNY3RoKulAp05F2Li+WrOTo4tTmdAAo
GxzbzpAdjMLD8bqaR6mrnYjFjmghkp8/DmpRv9sL665OSuzTXjIWPT0Ed24ebOQflxLA9Xfp8GK2
ArKcNBKGAVdnTmbyBoEBPOn0PEY708JsZ4oDEgObsRH10bFl0PXdDYmXy5/XmFFy+sF2Dv+3wtWd
wwI2zS8VJbK+lf4QxFZ+zv9pHimwQTJTO641dNyWX0BFmhTxlRnrgeWj8IoVfoV8iNrArM03BNWb
3zyR5Xv9Ie8Ke5S+h37Rks7nU13pgaQfz9JQacqVk0Qw6WXSPTzeJU5WC8traEO4IPwT0orzjgRI
Re8OBfWEtahPuST+EiadX++3JgihhYGMo8Kvlwq9gPTRMnlOu8O6ZKthhCBe3eCNwFh9FLyezCMU
nYdiIyIq/COmWaRqbqeNXBo0QyXf7/MlJf2YeM2R5sU1ZLCNzNqS8ntAVunrnBXId9OwGJEZeUQL
PCq3yh6RBwpdBQsGRvskXkEUL9ne3rCk5rmhjgwXzjTcwIUSq06YQ1sWdFqXXPqoKpgoqamoKRxH
PIbpua3c41JGe+LGhMjC4BrwG5lIidaGgjkuzWu2mnpGZ4o6tfeFQcr/OGLbJn8WTYpVZxHPptoQ
AUoF+CDFgqD82PQeVjIBbL83+kCeJiV8mbY/0v8RVtiu7ZRGZf+YiMr9kchjnLnWQf/B6BWuYi9e
BQ7Xyc7cj8dxfephg4qyZPDGl0P+cJYItvQVvcNeKmDgHyYesgfeX/uws4EbAUpq6vh9ktAicDBp
qXwcNkeqJD7WBORmm+3JS3IViNWSDA6Q1BvTMPVS2+L4M0IljMpHbWn/35PhP0MV73Bf1EiQUHaZ
YcKgJpkQWo8rO7W5tHBlsi441uZ9+PXWsByldeAxAbL6iSvxEKo/fgEMErctxqwE3Fp92C7auUyi
I5yZBWWXyBryds2qVMpxe3xggmKuCookDcwN2CZWe3v/X/8rsSK3sPtQ3pMdL92vXFE847hQ9iH/
LYT72Ms+Ak57xCj/CLXt/yFOqbZCdXBUSTiYurbrP8gRWrVMAfKQbFaeU6Vlogu9VBKvdTEKXV7z
oYkXMTBAbBLYG3GExbNGKR+tN7RS1+99+HX9/WXdqQN5amgixlYfqLURuSgye4IoH2SJHyFf98y4
g3bPby+pVg5x4vW2MDXDjbO4OhuxEQExBhcgRw2DpE5TXA0QWfQfeZR/XYp9m+CszqLq6vVNmyuO
U9z8NV/B7JmpNxYev/HHiAuogwbtx+lZ1NfXWetHH7H0sdVAGoJscA92YTTV/BUFlgOmi4qHEu/S
VnW1TA1kYHU1k9koKZ+k0hoi2hbA/Vw+D/OSbN6UlSbdvMa3MIjLsalP/oYwBJJ+/XiLT7kaTblE
wYkgUo+GlzD+BJ/mB+cZ0k0AyFZf+hokhQqqymL7YB9ZnACChRSpQ7IZVrMDZl3X09RLGWEILXqm
OCB/Pta1ri2di9n45kvWKpIu1oX//pbbamngPW6on3/HWcAJxPQbGyENBUezxna81KpiiYPj2r5Y
hg+Qs5Veyx2csCoEdmwpZ/bAniBJMxjgoYu5FTE2UQEwOB2jZ4Nxzp+GbUs55lw3rbtS24wayJfS
BGVQxPnQr31r8cqy7ivo4Wbqx4V7vgp0hyJQXdiSUmYoZ7AwJRcyYvjRji0Dru52mlwrHwsQywkp
t2p2VLnB7/RFkfYygrSCyumWM3W1XcGhCKL5nd7XEgQHdrPjPVFtO+8NNWyfynvdxLqMNhsnPoXq
6sRClTejqS2+k8wdX/avsQyE+e5P0G9eG52DlBw4YAz6QG+9u2r/Fjpy5/aTK0qleY2z1zWDY0pG
m89wrz+vr+N+LjqEy9en8hrKqQItMx0EW/yPHTY04kWUPMZsOjFn/0d9qgVR3VvjQuLuUtz7rES9
PGe9hyVMd3AMMSaLqhscHUYy9LO4i3dYS0v17sbDuLKFmoaxYXNzkPZdPiTS8INf5bfIkWQ5GL29
Yn0NSKy/EymYu6Wzm8PAZ30j3/q2Kht2jt7QnhMivzya++4OeMGTwFo2GNiBsMwgq0ZV2wMxxEyi
VpYFLu/kdgBeSJi7JMqFtFU2srVXCZzI9BzOxD975tVi02UUYjyV1ctweaRCHvVTx0JLt6Y27ix1
6WfhBH6EUMsWDNwgsXJ+77jD+fOO6fn4xck4DZ6Tr9bjquX8HZK7hdoWQRg+4/HQLk7g2HDyF+Jn
wYSqGEYmOPlm7kRvZ8Q1zBhMGCYpijU7pO+B0gpBlnjPb27Gu2BJd2b10PfSi985t4GxQI3o/yp7
3nnK1+CmjL5u9X+agO0PE9RRTNarLuUoyBEeBk6328VyFpYwxTUB3lMJOaeVGuFrFPUYzDu2x4E3
W6jmCHTE75Nwp1idp/QJzky9MH3EwvmFBQPlRFvrER15PrzkAgtFX8Jt7ng9NLrtwN2cuZ5H8Ij2
wiKgAh3ST+EQ2n93x4FiNpchd/zdYsWF2nnH+qA6PJ/LxgtSbIhPDwyIZa8CfVSEiRj7ALj03zLM
mDSLrCCCsK4DShCeBqAh0oO6CkzHIpn4A+g/LVVGkinsQ25ICRqj5o6QoPPfJB22QZFy3rU9h7gi
Hirf8zEOA6q5aYlcDXwrntdtxX/PqaTsKRSQ7QJwMsifs3hMJ+MgMi3/Fa51LsmmB4lI/oI+/R6G
MIUWWkk00vHTRGTE+sxO0LwiFGojMhQvirGmxoMI1QdxJmHPfThXC1jbbZ+tWtZDZir9hGK66cXu
v5hEL7ZMN9dtY6d8Rx/FMFA+hnL619exQr/aESOkGCf+2o/G5iZ5kz/YhT3iOPklTJr69mx6wHV8
TS6SNvW5IE3VsBaU0IcgwHP9vmj6ejbbwE9p3teMJIxYWaxkBb1nchxafk9ToqpCO9S2JfU9HP/Q
p4ulQHThP0uNDOLcYv3sc2sRijy5mHfdlslxdcZCWk1S2H+NIBEPgFj4p81Q5aOa+k9BSaLeliRt
85Acetuh/bWMEAzo7VDHAV/CAV7xNCrFGv+/Z+nGRrgTXxyAwxjzW0miMic0mp8/anoW8n256/v1
vvy4N+yy+aXa7mRMb8jcuj8fXj/y3D0gQ2yYSzUyX5LQYIWKBSrKq///zaPcejVVySKXhzPP7oWb
bTO6xKTUKipr/4Jl5SP4UcKYUioXfsjpD7Cov1kPn6mwWPEhZbPab+DmOVPqkLbmnjJlWTYUytGn
g1fKV18BU8/D8XD5bVYvPkixGjrlkzKRMm0+LrDqOOyM/p0882nhFMIKmEgaLuVR8ukj8HKd9264
32pVDioOh7Y8UNRTNgkd4aMxADxecw+ZjvDlzR5bB/BQoOtR+U1rJwB9mqsK9SSyDtfxxksebIEh
PPK95s4ekih1b1a6gDGa5givc4V2jv8AvZz6KxJSf/sK8tSw8EMbuK041KWFWKrv3zSk1fUIvprc
jI//57kqrjgEsE+nHIF5y3WBmIi6BlYKeFdSbLSigo/+dWTb6kzBd8cHtvzTWUPmoaeAwbkuwhL9
LMGITHgruCGkHAIFMM1XZeaVkKlTmj5V+eWyXFEfAjFUe6tnojb0LpbghP/x9PhAZ+lfdg9K+TCB
D5nbGyM0i/GVW6gzqm209AnqqkDYhKiLQX9OssDFov6gXtHWn1QHCYuJdCx+lHOQVISTR70CEwic
/xzFHMGeScCV586zeO50qJ2zVW4LTI5oGaT0DC7ThWr6UsgmLhv0656DsjBoN4HhZZ9Qtp1GqkZj
+Hb2YWVKAUwLoc0fd/msAsv61f09KzdD41RSkwUqgPhVtdp1t7r8vDWYh0pQJxlTLzpgay7djWgM
yCnefCLYSrRA9fdPoxEoaJHQMTxEmtSV3zqyPyrCo2yanzxmuz66SlbsWiun2hmEBlNdlAW1zWSB
CDbreoTGy87HUmwhrHbqZdmfUK7wh6vhfCC33epY0Lm2QPQkxbYD4WGVi35ttZMsst50m1JoxlWM
sbhKOTbjX+DEePUUNrokK9HnGXI3hZgvxcWQwwgLHzYk62DJ3zdmGmQQdsnI6Q0BRZ+oRnD5D3vF
MRj2nVEiVSm6vcF+/YUcgKmon3U9g3hgCdWvi9urSGiqQGVnqzxus06c8PErxzy5nS6CPb3oD+Cp
Y3+vg4wnCy85dVatSGHXaGCYbVUDTBgZTGvNlnpI0mOoHnHvPB5lmt8J5FhYlPbY8TYkfu0xCdb0
vn/nl439EOdMA8hXKssh82lq6t5Mx8iC4HpfZkFup3WyW+7JKDkq14CaDmTtV/3c9hbEdMuSrNm8
WcoZC3XkxgE1oEuO61bJ7duLVYLArL3o9RiT7NihXgxmJVAbXcGd7QSryhyOXQFpkqgx0hdKcCwG
rQmS9bUd1ygudgaJ66RQYkcbm3YMqBwgCG1XiGVxKFHXKcYdNXoC3jAeo2zhanbi8TMLI0TckvcK
K/ozvOp6dHqrClfVRMCtv/JngFv25y6+RN15wHWHLq3VIHkT+9Dzbt8vHvrv0ExgP2zSEUljPfHC
skMBt3NfuQzbaBowpMDkb0TXgIwRZjxIpq2ftnkmkXiPycZu4pV++K8H9IqykYLkGS2IRcZUXq9J
gC68L6oGho1scPPZDv1g505XJgnPIdELANjMY7Ohga2Lk/PolG/JDUwOx6+AXzV1AUXQwgZCTJMU
llYSRyQ6TSZ5EQ5wLdy12rcPJge5HLxh3H/h0vbAVG8qnbvQxhwE1dIBiM9y9WSJZ5iS1Z6TlInB
haZRUQAquX/Wm/9DSlLnDXpRULfjd7T3exJECsxtXNdxrzhDlM92Kyj89dIawdOk8U/qsFVQ8K05
Ufx++Kcy/Kt25Gjg/TRxdTbWTdSVLwm+ig/srhJeP5ueF3xiHQ1/rCQm1k5LZkIehAxyDuWQB114
M8wqJY1EIeL4oWr7ea/KxVLto+XX2lA/dwvQLzxQ/6eEzY+W+e9pVA8QObNxZE4+72SeTCymvWyV
mp6uHLY/v1q2MHyxdMIOzzaPjlGIU0xuAH5TBPy6R2n5jMK/pV2hHUVTojAKVOsSGf7kK6W1skR2
gBqVzt9vCoDdk/ko/yhwgg9OjEyBRYWX0ILozNEtBG47Zs4Tx2UBgJuS7fwti4dmvInYJzpfgA1F
InWLyDuKAcNGXa46J2wIKLxjFNMK3PhNySsmvfPC+e03iXacqEWzhIXeHKY0jUVwZEKhyX7BVLza
xK/frwSDaXFFbX4UQdgx36rYqCrXMnQxUpWJwBawQXYoMW8yMTg9wIE8AvDi9+SZ2PI2iSLL8wh+
D9Dj3jKRjndzM8O1Y1CVfYAqlBpL2T83fR3ftQEarQ7ZL/DwZHnOPr9K0uw53Oo8r7JnTrLMDIGY
WOZt56eUYXhMGqzAw99JSXoi24+51X+fBa+sJvzRMIeurBF2hvXgf1jY6vp85xYNTOFOaYQ2RD6Y
VTWL081L5p5GeaiDltc7WbfF4iQXy8shkX2sZkunNcLk3v8ig+bSzV6y00wvaX+b29IpRQ5IbaWz
Kofo8y2rJ1DQwKiOcfFbVARPu3StgaD0NkjTec5H2jXsjbxhXNQInQXlNA2Y3yT24cMzWKAlpHCR
eAgFj3RnknRsDYzSXXvNyqPt5jq40V/rxPyAt5NVZBiCh8lBVXoy/UlMxYA8ufX7YuJOFB9gQidG
KTUKi/R8dGQKHjYzGhPooIRdtqnI1KhnrV+R5udMJMYVdG1qfNDDcJh6VW7Hh4mMGWs7q0/iKymk
1WV2Dxi64E07FZfJ1kCfZp+hi/c+I7bgnOihDLCiPS6QR5sB6yP84xDsZ6QY/ee2iwwiumMbGi+9
Kr6f7taLQ1almkOsMEWNtTGaPpZdtAM56sjH/2eh8TaOycvaBMHPI5JVwW4Bv5+r5Z0Ge8QbVHZj
VFG63CARV1VzJkyX0xzgpH4pW3BwOOEBevDI3/Ik8kF+oZjXjAyyUOi1qGuoFHaY7EpHsxI1xBiH
Upsy3byXSjvHEvbjDE8MKZuOv1bSde2rSHhbi/DE2P8zRTiGCKpTKKAV26zAQ5PKpibWi3qbXQbB
HjxMWH1QXis+SZFZWgFfGORh3tQKOjT4ExyXJdUTX3Rm/sMEDZhJgdo6SJfkCYs90Hr6h4wFLIGB
zpF4YOnPzerQfKCnD1kxAWMANaD3E8t1qAKYat9E/fRWnVVRf0OUHKlR/ubYSaf6TEbR7mHai4ed
zjZjRZtznlEdSOvg0HoojGiWSrM5qwra4Ruqk9HCiZM7Qr8FttQfebqCBndlakKzMvq35Jb3I7mm
EcOuGrS/6R820ma6c4hVxKZAt93pnsCBx/uevrT9a97vAzTi04HvYPTORw2OBwh6aNUujR1aPYkU
7cYDKoEaVJ5UaGQrkiFd8dTDGf848G4O1bpooS9mzntaBBL09s8zssPamQbxMXFdj2vcxh1pxDUT
cDSnsNp8+gxXqvjusNJ3EfMQbpceVqd0Itsencll40g1FzKJ83YPm9V8x5kBTM5BWD03bJNd9C2N
1lW0vYbGh15s/f7x0c5gZjrxXigCbEtV84RevZFMzMe9J8qVvtRkAPg7nlg4ByfHNgOkjwT3mGsc
78a1fNki2En61bU2BSSwJcyGXjvO6da3NRltMPc1IBJf79Z+DsIT4YKECowF/aH6DNbIaG4A3+Yv
CjeHolBKKRgQUkddN8iVndcEWhJ9OidIcfNUygUNSyPFPnewEv+syq3aCVhWPzi/SX31BqlSuI2W
rFyecErWX0xSbMDFoRmlRUsQTT+jc3TGkiFPzvRrrB+3XCqPU3qYszidySlUPzlVz11xD2kOwnhG
zIDpauFNexFmqJclNFc+nzOakjZJVRCpysh1dsoXj827+5ICAIGMoYNz8cvwKLIlmA8q8Qlgf1Yc
d5UsSyWV/FYgTsR9nLjN5gVFClGu2OXbPOfIIxp4VQ6FezdE1OTt7Ai25zvep2txF4xuYZ+zDWEb
Z8sG2O7fxfe3NLGq18zxEYfrXBzart/xK9g1ygfQ+ECTCCr/iOMr/BIUfB1HNfF7E2fk7A7D/J16
ixzd01YUhF2XdAxXtoi4FQKheArdBIJpRSy90q36cyzNs3DfIMPbAWePFgF8T8qbsi745TVpBbC5
IWLYi0hsdp4EwaGQi9xOsEQnGt6iB7By/K66dRKTHVr6fmC2nqBAaQGTB86TF8WyqOfqo7UoN+xe
OSOhnbSbdoIiuleFNjriA5SvALgR2v7TfQ5DXSPo50WCE2br30AKXbp7lgdSzYKkfexeOhFpMXfK
DXr/lNalvVoeNoUgIqn+VhCp+Jb8NVhBCEKsCYeyqZkziEcccXjDhsvovF0JixnVv6EpkMiJWIL8
mCZ+SEi9DuP7UqslRD3ehAqH0PaPTDxmsLf0dsOY7bqnGYhNNy+H8WYStFoQDEihvVhuCdfzVoVQ
eGSGVyraH7NbR6bZCPPQC1Dk7OigvftVYWGBoX0ARC3QO/d/v5d7eQOIpJHLmE6lxGhNjCN025HC
/lriI61mxzUs4gyQaFlQJKxt+HDo85VaJPICTm2IAalXc3HBjy0i0N3MCvFPdV2BkHRjDZUaE9zx
bGN0ztDed+LarWNSXvE85IWb7HoclA+cIspIY48mg1ospqNdrQnZHLxJq0sOUfSygx4Ybp52RHaY
uNO7i+zVe2mrDS99Fj/dQpylSMTF4h6IEq3xwPCMY6Byh0JBQNdwuBtl/lOPTSD25zHphoPv8Jua
vBh5Tvb9Ji87wtIN9Op2WEybdkUZWlcNF7PHTdJBnI9eCOeot7nwxzP4ifVyNOF6jHhR2XCTkFiO
UCen1b+67BciXx+L2KSFUK5ddRgRdvx5Xvl25rcWc/P52SQ8165R2IZPgruk8DXFXuTWWF7o/Ljx
ZiPccLAERfHxTRLnoLGcCu8RLPpNhUo3E5AeI/AWx1FZjmkwNchsEoDPm/LoZ3Nya8bQHlhn86wU
UmNz/NUoSj5GB/rPNDGdwX60RL0hcSoY5QhernZb/Euw9Lb8r5g+crUsiuV52jH9z35ZYFU0xXrM
EezVDheoU91fSTZ100peU1PjYi7uoZLlxOdmjnJ+R41soZSfhKjFKAXX9jNWITVdBPCouiS1Qov8
eMU9U3K1OvutCxrVIlJOkWrxyyGea+Md80Zh/n+nW21pVqurXAOQEIpc6JX8m6x+a/ttc8mZ6fU5
NYIYAdYKt6c+F5BYRdAwenyux6A4afsZu6aTHWcR0QLuIMTOTtRcrknQi6X/sduJZs1Sy1wr2uiD
96ZbhXHzBhz+0mchAQsN4L9I9pzZ/lemR588LDUQwMOoEoQzsP6f6Q9GNz2uN2hizhOxV3c2LlzT
iX+i+3sBkV+RuuAnPOgix6F4eKET1U2X1FNuf/4X2rtosCgm9G6+lIkhtDjQKXufS0hdFIyf2oat
5NxsWuJnuYuGXLbcAgUApiWXg7LE7WZArsZrwTEKe/flWtmJrYcP7T9/ZkmvIFkXuDQKb4cZXSDM
ZzY2MBSlnPAc3DlMu/Q6HK6cYyNAKT9AawOQfEoZywGXtRaw6rc7QMnt1WGEiK3ebP/aOmQ/uL7v
Obn28cOc0/BJXjUfJxwW6H2KUgRhU2kpQyihk5K8/JqJrZ5tG8nLTip4nMCFSiXXjCvJCTIfBQqf
l90LSFCQYqFdcjMMsdLxBgajoBlWISdDoSSkmbg2KAE0D+H0qaNYSIIFKPu2z8IdX4XnONNojgkP
ieKICpqfUt1W1QXZJc8a8K6zts7begQZIVBEIYL8lvu9Mh6mboaiTQ9pC0iMACZJRkYodrR5CO6F
WucGsbyIvyaKZBMxN3Yjj7xpc1XpKWmoc2JHXC4hAGw2LUrG5hRgY5hV/CT6o5VPYzr77UvlT0mz
aOJqaSGueF/80lTKzZjwHSxl/A/rNeCYe29LPJE0Whleyd8owYVRXmWJ12Gvo9gtmMltvbnwAACA
Ukgx7paldDOwxjFuqV+TBvMgIj6hMLfx03JEpR65R1JpYEnuulrqPI3pgUXJDftGrGRfELH5z8i7
82rG5XyE6bbm0qMLmpPnunCv8TJzcyeygetaZ8XmZlZm6YZLVulYk2FNjk4S9omkrjj+A3jZzAWJ
rMK01FvYFRLW5hEK7VG7wW6lf8mBnDwSyYbBmqXGi9Nln1x3CdWAfckGSOYk0mElQxgva/D6uZ/w
o0K7JGNf6kNfO05isJtJRjWay0AYRV0fw3sOli4xQPqe1c1JFoCXQg0F3JJK0jpEas2vohnpxZun
wCeTN9r5rhQygyevSkQy8oSkU/A9Kfdx2D5midO1U9zhKPf0fdzaq7eOoCaNlEOdIKt3vcTCGmr8
ikHZjGDJZlPnvRMVmr5sqPLDm8Z/EYh4pRdngWYNuzOZn7+N01lIkwjat37jYHrMuxtr16WlbpFZ
KmAzuGB5C/u1ChCImj3lbR2eC6k0kpmYgnANTPDIkzSM50+bcSn3zA4afoBmysm+0xORgagEiiVG
gVHCx4XjfpJQHKI9/VicPaSM+c/ggnj33nvWSCj3/Mxr2ruobpmb1T4F5C1gBEAKEEX4wqhtSQKd
XKkUF67s8Su8rM6vXYjGP+2dht0JNhL869QEP42e8Q0IxPlBkzVN39WFNsVp/5HahSkj9b6hdV0B
ijaO2QBc2vcNyVe74qSebEMHSTvEb6MiUAdJdLoFWL+5OoAWs/pQVPQcwVER5v9173to9NUbtl1v
w8hjOyTXJ6m1Okjvu6GGvR0jJYnmi8Qr7F3MbGmn392t8dhH91WkU4W2wOaRmR3rditksjGzcgmq
oRYR8TDxGPSqxSArA41lpUHJJCcOQCbp9e8wahzpFpaDCNjkjrVkBRp6horHHxWPGL9KrwRsl+cQ
0FPPemdrjIdljKW78fbn07VvnDi4XiOXJB3qbQqxTpAGj3+Aw43wwL809fF/8K8m1wnoRKYyfPvs
x/PJz5S/GPWa5Qvd/1Bi11Na/oHfusVQ2pbrd4T1NhD2yqNzX4au/ACoch187mnp2Sx38ABW9ZB9
4UXrCprRgd3u7hywIqw+R2KKgQ02emS4lVK5PKUD/f8tSSLLlmd9n6Y8Z4O5TgS3YUZRHUVbYL9b
NlEyftXJJ2mXICJ6d8CJJjalF2IH1niEqOKCzXcvmKXz9ORNTJAc61B2ciVF12i6jF+8nK4cAMQ+
x0Rhn9KIxTh27UKTVfj17AvXiq5qbsbghEKMuGrNqc4z23VDEhvLh8OJq3HG9U0ga/j2vupu8AJL
RxsT/IyMYl1ZUiZMRKzQUat0Qh7RLsXoyuB81pTxmJb8NpcqPc1HSSdFZj67BDnuQ18/plvn7rjl
OglUJOnMBq+Ovf15yOgC+hazizYEgFs+7SYEqG9oViVDXDDnWSKOoZgWo/CDYZrHpHpfHXYevRXs
BdMNiNQhVWP1u+pYAh8ZiQJw5BZaduCLsolLk4gyhrUNY3kwxom1JQJVYL5pK9GY9nxa5bbUmSs/
GcGjswGM7BNu8h8wk7jyr7sabQweOr3RzUpHCJMEvNTUUwv4m0FNG1w7of7NewYgQnXf9pvGy1fJ
TLD3zjW8ONuLiVnWW6Ia19eLFVeXFZB9dRojS5U3TdJRR5GNO3X6TL4mnGlVh6Im0Yv79bnr8dmo
Z5+mp0X+VIyZiidUocWFtWKg5OyuVf3ujdsqPlXP8/FdLoeGs63n36CY4/E3ZTVLt9JLpqQgOq8O
B3nqclJqnIu+c7NZXz5CnSMv1cdM/aboS4i9Mws4pNrUBlqmtefwQmXwxOr/Dje5Kd6amGBnpVFi
tpnoFxfj987Y6Z4vkmf6h+JlmUag7jaXpFbakCROeRLUYEhekb1h2leJamYx4idv7Kd2WogBtSkg
g7pVyTtEowkForGsNwJ+mdlSWCkC7mGoBH3jGa1Waxq0PCsboCbwQRxwL+noPZm/jIhscfIPooxJ
CBW9HP5leh+AN2GJ+FXwsTy1Zd4jWypLe20+sf+j26KSVHNmu4cIVnV0CmvEs6v8zF6Rz2PB/Bfq
tfx95Rnfhq2Di13jCF5GzeJ531UgtOAoNCiEg54h/D9oxeDKuU+AXs8+CsEtTJ5EhkKqVy8FuSur
V41Dk9u5wg+HbVBJ7HHI55gmCpJ1CVA8Empz6x/KspWgzxvG7NV3v1c5y4TyRn7ruNy5ecRensUX
U1kbux1bejuDsXYvk7tZC5j+HAK0KbW+PAtu+uWrGw9bO2e5sU9Jbpmi5E++KjqcxTb8o6IZ80Ci
ZRqwb9s2O85h9wxWt3TklJD19L9xe2OoYoHuEXkQq80+cc4eGjwyH4icujLqurt5sttvYqcj+sLH
zDuzrW391mnL5kyC66VBw+6A2wasgC7bXHc/izwdGtjwmhXBm6khA0oOxZllo83yE4dKsV2TeqWK
OzcWDlU4EdAqpge+2Bh8O8QoM8MZVczVtzEGD/7FyENDuRKnZzBnwKm8NlC6IDsy6V998LeiTNlF
V0XcVjitZk/vU3UOgaK2iVcv2B0/v9hMx3nf2l3b7z7yuYENX0Rx1qztfkb2ezaa8qzQCSOT8iy8
LerY1clwabNLTB8DTglhbOJbzOgdnNW6xqCENd9meD/sk1ekH0aaI2Nu9Sof9dgmFkt7NRvCWIdf
KmWwwxkHSlrJgUOm/X0P7ci39LQaoZ+xctHjj6n1syQC79RDFYXDgHvu8YS0dqP8MRvZHKoykK7B
SA0CfjWBKRBeCsrYWREPEpT7zz/sdyOXSQhnSjbTnuqUUKzeYemdib7FRiEO24v4PvgU8/gTbqt8
E9IyBHAksyCl+MwCQYyosimRDVeAXGbUPgprjpE9t2TSQFvxm3wEhGONiEmimGkWd6wn/NjtG43B
RO2bWGwOm2nR0+YdXs0/M7wkBhQATp/LU5ClmM6aTmyDmRqY/l0nXK3loq7vIsJQHNZMAH6CyCGo
TYh20m9v9k6NPhmoobZ1sJqAgazuSHNI0MS6cleN0AOGMl3cqtWhOKuVFcYvq0Qf64yEoui5YQ/+
DuaKHTlbfPzRVChTQEZ3UpXepto2+09S/hpVaEkRlbfSd8Om5BEjRr8GkxzgEn4LuPvQv1Ld/6Mk
L1mZ1XkuCYN9xEsusBd/uulLJ7BF3lFqritGS4IYYY1Aa8zm3sClLYS2PfuqMLEw7kCJGajgAScw
fNMMHa58OOCBK26JYfWgwAKbAH2MAKNrXicZzx7VeU04KHLxs/W/h5zBV7fMmgD9OCdhktvx6eaK
nOqltSMSMgAMv9tSoeBF0Rr2A5UNhrLOpp342vW5B6JLXQFfwSZKtvjwwGMjVG7FABIc1DhIGJTp
sZeK+n504o05AqSCWMtFZ9doD7jQt3PIDdcDb+fXGEHHxrK6FY5hlYdqLEkBO66WPoTAb0Lko9Xr
oxjfEfXe9e+rY7RxGP/scYE/lMuLKEDln67NMpH/RLmVAezbp5P+K5ranFpYpYi8ya9YnL9LmJlJ
7VB/Do8OX4kFCUR3S0HXofLHmtsSismYrk+xqkYVOXnbOzadzaEhqxsHn6v3jK99k1VN83wolHZH
M+4EKhRBxRZT4fxMQCQsOChBwvgmTBRiifEMkmMXJFwLvpihEOf4XRCnSjQ8DrzrZTps/QC07tiO
5wkX48YqBB0LIcX+cd4FmcJb5UlzTdJOKbz//DLDFO92LTbZDNZLOjKEfGy2gZCd6wMi6TzU8Js1
uDIK9a8UEgTozV566pz+5Bc9DJ/sZrz5h1PkyK8Pj9ZEFbCLDZ9pUYdOBnoY1H+d8WcaMQS1psC4
I12EsbTQTyzJ4dWht/61V+9pTMJPHLeHAYySG5tcp7OIw6nMkL4IPTusvckYviDBeHyMEyB/sCkX
bsdClgXmumxNjbUiCLmsayyNNCW7sA2xrzwNhgkg2RpaUn4pouEse5SgctuURfLfGaoXuHTTsdRs
h+F4nJcqLZi8Hy7HurMtwUf0hDkfvbE48TBcMpgAEETmV8AgUrKCnCrEv+dx0CzDTvOpgngo3XES
1JX7Jm0HQUB5k3rLtATKl0+1EyR275Q81G7VxkZ3fmrWx2Ri+wowCQcIiqvo3cqvGcSLgQePjYyG
dTBlqjyeurBBKxetavl9AjQ0J7/I2TzDe96wkRKl/YwGu+ynEOFNh6RpL1sZG27n37kjfWfqCjL/
P9pXy/K4x/dDfl5JrJ72z0Q49UTY8Lfrj4WjmriEZqOW2RWlnLtSWQuN0DJdWPwWMMJGZ7XPpq/+
mhBGn2HmQihffiQqV40j6uo8Fl+n63yULKdjRtDDEJeg6qNj5TTYj/BQe8H1UowTi6afvu0d8xS8
3Y3kuWNiC3ZsK9UkihVT+FdVhXCxPvoXMxkqG4YOfreA4llb3J2qVAMI/7LGuqIdZjOVdEVnwzhw
0rten0p5JDWE2WDBLsQXSvKWcCSHdQeR/QDtul/geg8pEYSVkLjmfUCjXV4wvKnMy0YOcVHhuS6T
Ir4O22iF84MmJ8TaXRKjVjsNfDfdxI56u+C3yahAKTTJB//f3LCT/d3L00BPMGY0i3L37ZJ4YI7p
y4vd0HhtF/RrOpJ/G1qWDIspH5pYm5BwXoOi30VZVTBq2c7Ts9u13sJetvKIRGA1Sg8mn5gd0iyC
mg/G1eQTdWVp5lBq1YSHSVq3girEaJ8MKuaQNYjuidF9/EXBD5F7fyFmqQf5zDOzBlBj17Owhs26
bQPFq+5hUvtfCaYXZrRkfJU6hAIMafvgvH3ElU/I1sQEPvZvxPuIr/3RFFxZog3hjedY/n2e9VIH
v1WZx1CLA/SKnGK5gr9CRksZdV07fFofWIoViDPVRGLhNx3sz80+Qy74ubsBEhDlzMUw8sKZes+U
Sp0u0QNdWYZmLPtJk9vJoFdaHxyiRHeAiQS3ju90iD8pAsAAen2+NEaqs1OskC8HE+cIORzzcS3y
JziGgDg2zIVwKWLrAC6M71onjATLsQbkCJIIQ6SPvAjMzinVblO3WBQK3kHigVNHKgd0VPmpF2Ej
6hEZ3L5A000+ffhp0E7TKUc8cw/4UTmv4/KCh27lTlk2kruH13uvu4u+BUXhafNp75Jl6TbyW0R7
fPgbxmS9naDwuarRlqJYq9IkNAec9l0bUod8inWGzR2jdLUql2wZWG7dbivTfSdj0pmerbS3HL8R
cgVot/TSD3TiRBh15uW/nZFMHsuLG8QVMA2XTKcU9RfMxUYgb9VvlKcQfVQUleczr52hNwjapodi
FTYKSYchi2MaSv7bjcE+Qh2IERPCq0tp5HRSzh2bsxsEnK3EgklhoYg3cayl9khROUO/aM/OR3dF
mUGIR1LKl1/WMrlRB50wvsDTCs+x4mlPa4xRwy0sV9FoQx7xlR3fNoXGSzK01x3SIHcdf6zGfbLH
Cfq+UnQdlsRXFOGcuUnv6YM40VxH9MZL6WUPXM32KyhnOt8XF94XiyqyKTvp8G/t2HCsRxjAyfxT
txIuQ+qHGnRvDMaEI9YYHV/TmkQXevIty1/5HjOYkcVXzzC7WtuyUfht9N9kt1q2fvJMjV9WHap8
meWLAtomjXHkWrJ8XpdWFT6WlbEHqhjmX4oyY5d67CqIaHMKcUdqD6+0kiF7Z3FXGTT497nMLDnP
rURopFhjDKQaN4yd2LP1xdEPeBET9btMaGDU6UiDDHnRNRRI2HW3tb910ghYr5+IgjSHxZAzNtk2
NSyw8YtFBI/eT0skaiAri9SUNyXnviXuNzG6GNJsVxFLCL4byNBHSdxniV2zATguROBm5ylvf7+8
qIqIjrW+j6ye22lHJh3g/ny2MVsyZoVzAEhixE5JHtj08kEK9y3BK/Yxv2IbJrE3mrVqV/rdlBiG
X0pDo8z+AQu6sVZgMrg3Zj569z6dNhlLVHbXfEa0gs7L1hbhs+wltxBT9wf6YTSyZsOcLjtPE675
DSRj84kwXxAdJUchJYDzPgKX0x/rGdwqjUti48XZUPHLN9QURKaz9IasThfXuczzvwfcwZCT1pS7
eyKrbXgyl5UQWIwByRAAbPtVtbf1ZTw99BH748acS6kHQLgq4ltSutBv/aiGiZlIbkiejV1KTKmk
Gy0iPLmUzSAJPT9hv9e+gN54suD60jGqIX2GmsRuLfia4TsnDfNGuDTj1y8Es7UwibXYLvpAFZfV
+70c/avgHZ+k7eURpogYInDJF+sptc2FN2NepHcGdUizT6ZWKj2QxoAtwgq3TTYFZyFmXGFc1o3M
nUpsxM3UIW4/2QSZbG/fukKPMefCX69r3/BJgTGS/cKrpL2bZVWcuIIRJtcJogTN0LndVQc6gHJ6
1zIxfx/Rfje/oRx0/pwyazn0rq6u/xxj3v6e5IM5+v90AecLCzHP66/SDB6sVhxedNt+D7jbtFSp
ULhvtzoMrUyiQfSoDyIUgxFjN98lKOcgGsLsDWtiDJRAISkq8txQfuo0TuWJHt9Df8DpJ28jqwmN
yx39uvAsVzz4ZF1joWkLBd9s3XeqACpkP8jlCXJziF4ArTlN7NNbzkcoZjGeb9OYeANvRzqQPgJB
57THDzeiQv+GlA0snFccNgm98H1cUHPS3HlENM9CCovqnNj/EJ7ehEFcQuwjIz+9UC+reFW8FPEq
KBgpqMHO3fdr5KmjQ5/NEiDvaLh8CJM3Mp54PFkXgtpMiV6GFwQk8oAdaxaqJ6LSOFH5+cG9SvaY
YQUoGvKceTjDG4Y/d8pIIaCWLes0MCO7S7FJzgQn6/WBuZ0/OPzk9FJtcRSJ2vCipXzQICW5VNgp
OvVvVN8vJa15pQs62pTG4rT/a3a8/rpAUQO7/jE497jiy3zueA+tc4ZiiRFbyt9S1SZt5GmMtWs0
sqozlUXkMeC6QGC+0e9H50V4gQQvFaLr2/yZuXSet/qaY9bMoNdAbZRelf+CLJreEZ0m6bwEepB9
OvcP5z6UA4XANB9HVVkqT+JXFdvLTii6O7+5cFk5oM96Sl/405DxspOJPoR7K30dr5KrTjc/vzT5
Awt4xg6CcJlK4yxHS/6MXx0c+pycbTTaSLa198/Avj9jUORlJUDM5v6TH//LKjU8hPIUi5pflFJI
WopDap3gz7BEVNMbGhEtf0q946zttDJTQ9+5xFyZRrROqm8IXW0v7QJjUJVcqekEJ56dNaJckqnz
xht/lSsxVEGPespC0or1k+MjsMjcihcq8VMMGd+jTcrnEfMryry+aN3Bg9LtulQufxCfWGgQ7JNH
G66+Fa0u9eW4Guu39CPRi0Bl+UGgEXHr6BxCXNb6KlZZeQ4l6sTyeXAEtd79hsLXEk/22LPXHLLe
YdWdU8aFjojAQEOqGDjVMoaHkW93f6rEN9scMmbdPIe4CLaAhWBBlkGyt+/tzsfeyxtUszdZxhHA
fEFuCe8AmV2T2cm34dsDZ2zz6TPj9qbFbhUoiaB57Zzt1xGAWPGApRI7q0HySA1zuPDiJVhrx5eA
yvcuUatLAeY8UuJOvkDK6dovScvWXI+tlP/A4sUUyns0kXpeh8FuiQI4Z37YpbRHhaitdj5YWjTw
e0wNAZB0gVAC3hFV+4FS1217ZJpM7YTA3LTtlVJ6bAu3iNdXFGPfJnt/kNvoRkWSTjEyzwRh6pNi
7w8cWnx7xDaWIEVRbLB3iLX8PYFxE+w5Fjz+hbE030cjdLHbdG9e6G4SXXUwF6s+RIaMNjEC/euR
F92zUfE0NYBJ6Twg9grIFgxNo4nJTYPQFdbDGWhNqUITee49oNUMfggH8ph4z5fqATU/6HGd6AGr
jEVIU5dghT/UIqVNw/+Nvjgvggrcn0YuE3HSXm7+bVa57va2kiAXRRMHhlQ5Ql2dPquCBbf3t59V
WoKcIXzuNm3fhAuDZpCQeHdZ00CyD6On1ae2E230dDiDNYXdmLRoQOpl5HPEW/cGxAsjz8LEiLNq
SP3xtKo4unkIyyPxF2b+0XZ7b0VqHx0QVLyAZrPNZDIYbHRkyl9IcA8zutXmCQewiDZ6LfgbxFpZ
dsaKXzOG6tYoiz+lGIXJDPfMP59rorVg33JSGi+BIW7qMYabJdwu3rMp8fmnow482z8FEYDeRNpT
8PqMaXmpT/yK8xDVWvU2gdBMYsSR2h8RESkclscyT/pqCKaL23eyC8GPV/YupnooHO/qgT5azvMo
JcpfoVY2EER14g+pvJ/Ongc9RoCeVnz8909dmsNzLLx2r17gvPCSU3I7Zlo8KqlvtTviI22UtcKi
2IKIGlqOQyrLty9iAl0VAe3bOEs30fRsmAG+SlxFNpdfrXThFu9CrmFuZi0BX6xjOqTqWEegqoaK
dL9Xgu+CnUX4oST/TxZH7ewygI14Y3W3t3bXkRLQXjGGYLvfu34Dz9FUAyoRhnMtzwnCOEkgcT69
lNHW7kprxmzeNI4eGwSbzesffnPShml34uKF8zUzEcL4qe6Llfu/Da+Hkzcq3J4EuUmftK9BAEvM
b9BmU0R4wNWvRpaKpCtDbV2uGmWWemGn2TfRTIBgEZ+iqJosGd3eYhwZGGbKSCm9ezibzMKbQM88
0igRwloZj7gT9rU4ZhA3tnXGmnRtK6l4rmWKRhFm56Xg0viaTyX31ZQBCXUVflaPJl84SLBj/JM5
POnq0JJYuMOlFohMqmNe0Dl83niAiu3xw/mQM6AOf9ZTi7lnmsnt6wViJlOQkDJoUxSi+2XYGX6q
1CFIR3x1TRMn9Y7Id15N6jMY6ogsNp8AFYd3AlvM8xuZqOVT0huXucULx5Va0sDeYzsaX+94XEp/
V7v5Dzmns8NWa4NWtnPkknydAZj3xJxy0SafDw9tfenqlE5YF/23UGbAYR1Ceuddn4jBjsmdrhd/
doOe9QEn7RZp2516za1iQ0+hOVCYld9t2povhTalfRT1KJancBorqciXLGNrsOx8N7nFHyxt7j8Q
TKFKbgJRDoXCJ6KNMH0c5Y/7NQhlYKVxcT4k2dlXk6YU+oqUvfhY8y3c27Bmt8Xqcw2+ZWXis/yH
RiuZA0IyhHVCCPtD/ZxORu67E4qjomOylKaF6TQF14RGudR8HG9NXLwcqaxZPaiSd54fBxFDIRYA
NpzoL/zPgU+o0OndDOluh7ROVuOR8/5rnU13hVn0BGsSQ+NVl8tDzg0SiGjarcrkkyhmqiIWpwbS
+plP4lJBZL5xJdLuDjqmL0jqgf2wQfFylid7/KKcr0oj/rHMpIY6Q/tlIFqCQywBNSDLrcoE1nS3
DhqR/e9TsC+MJ5xe3fCpR6KG8dwYnxt9vIOHxzQAlw8Zn1BE2INywfn5DU6W2AgqwNPKgwbBPIav
CURheKGuGCWP/b9XWwJZtjYB7VkGU7mb6ZiZJR9VNpf388ygFj3bH9WOApcPnghjTw/DQ7TELgt2
MyFE/M4KwgvjtuhrTb1ep7P6OWNOS8Yi8iQDojw8nlrgz6JVIvO6mJESS6jzxNQf/bT6TMXuQPhd
5NDz8v5e9MQVuPCsXvSCjRGYO0mj55ZVhVmmgSIUuFKZBcnTmedghByLWIwZuJGaRnYWhKDIStTi
4SaJAajkfPNjLa3/iw2CPBYbfoXBqteLHUfmvvuY7tTL6nPQ7KFpT1OyjCOur0dVIiHhN/nY/hzl
uv7/qGigfrmKSkl2QJSM6IVPrD/OpRdbX2MlV+pEy9s+2K/Dju+JSny2P7EA6sJCwbDovQK46MVT
5aseabNnz89h7IF25164m5FH9cemD43fTGQCNXcvo4Wp+T7jSIFZ9vXKyLs94pIwoqTBSiRr073P
1IZlWr0nIpSVMqTZIHZ3gWHQ//E8xb05+Uq/iYTsic+zUu/8Px3BZMGi/o1vZ3xZAla/8hHXk+YL
Fgm0fmtOmi8gR1S7PzdPLbb1xRp3tfBStws8aYotpsqiIElNkx2VBEP/IFCVITRGfUj68AQNa08/
pQRvno3ZLeru8jUdbCiKAnLjhMWaQ0Zk2HBDCiVmaWRKI2nMYsJ+h7Mhur70n/hK9+4KUgi4wGzq
2t+J04e/ZEB38Zd/WG83+l5IG+6pwB5Vx8yKc1YiUG6pPB4DZELdJuzw7oqZpvtqEE89RhaSkW5Q
Q+mF8rRdwEwT5BU61C3dI20smcBA1zN35odnkcwA2n9nnqy402GCaixK2nLczNdXFmegBrdklwoy
KsN2kz3BGtfwTW50tndJI4iuB/bPGLcPyelHCM8UlQn5TwBD8YX9Sr8YUw6W00CWLtWTMKMubFYm
vNw0GCHjKKXPMsFz5YyMLew8Pgi7xzbkQHxVgZf9I4em0NhRav0/n8JIW2qU7eSCVjhXib0yh2/w
PmLaWIOeHAyOs0Nlay9v8AyTuFTT1kqWGS9UTYOBMLlWCk+BwnW9rUjRkzuC6E5dPN2wrC4FXjPU
gspaVKx0CC+iON9HPMSCfkBgrfM9KJXGXtK2hyINT/xAjCopY54U4YGGNKA5aM5UD5DUShq7Njs1
aCKdOu3tx6i9BRDZKPfW5iaUqZB7PuHW31odIjRlJj2CLdOGezPfxECC/th3nT3S2XphR2psOWUz
IFHFb5IOKmsceOKYMKqz8PYvDoH6xaFHLWkw3hCrF+VVIKl4RpcezoAfNKU+kBBMKig+NpY64vuO
Iblw+iylRc+RnDn3cZ91EoHP8ql6k+Ex3UdEzHBLh1X4NMAepKyFboCY3FI+M7J0rNW6YtkUL8cY
COF3IkPyOoGfp3wPgv7pkq+zpbhHUYDzdUGLGTZDANnOFVfVUrsrht6WzGZTTapISZK4hkmXuEiJ
X/IqH/FiF+TO0PDot8q8E6I/atOj8hY9VunxoRA6leV/apJVHZFymLMFht8i9THjftpu2oy1YTOU
P38yA4KsHmQYrPsNeYqGw6W3pv8VrtZ1IBGE4e4FUXASM0dWSWtpYdnDdzKqgZ25jkyklA1C0DzH
El7wA1TiE5KNsKwgFsneAwFfz6S+E5rae1uzaSzqCgxW7JGAbBFa/UgInH2kh59qkCBoYbRakhSz
lezY8ay8B7SpIoiuRQBC/MhGlpkw5oxu6vE8OF3+qW9YiBibC4vbxu/9PTz3nwbnh3TiFV+bzk0y
3qaGN5LOO0N4FdhO198mABXnZmjGASiD/bOQ758TcjUCMoHrHtn8pFcpdfu1z0duLvMuNHDGHJJg
an2IoBd/kLBEusxMfW6tz6S8YU4I6l/qEsE1tHGp6Mm8bnfBwzQz0p5l8l5GZ3tDDWPfgPP1Cd7u
pxPLhWDcv1qbqr7UBb/bwBfU7g16vqZ/3bImFDR3Lpevl/3PQLq6YET4NAvF36UyhQizAW91mloO
e04WkZurontg2dwO8Ag2StbXbmL+7DqjZQ3kNlqLZs3cTTXB2q7YJzfQX9Vo1NRHQOpbeSLm6Xzh
59aoh+uDoAzhozbQhxlox6nvUmRzpavW4WiRf+7SU99Uh9I9ugr8GcqxUff/rN8gta6SI/nmvLUN
M5dn9YUr2fKSDvg6udQCECD7/74lr5O1Oadnf0bF50oG8mf1g8/OlR1qWs3AFeMasSR5u0VKAaPg
Euu7BdxvkZ/VG4QkNqnrsYIsCdn1TSpWmNDWE05Kgqnva9PaIV/IU9bueHgVmOw3WpV9LtZLzE1A
gq3IvN069q6oN7t+gz3Ash9x6phMB+qe1ZLgMlhVi5xgL069AhNZQRlnXoE82J8Xbi0rPtJD/boU
l2XNABl4F/vVVb8h4KNNMPdA9SxWZRm43Irzvxp6mdNkydrJUpGEat1vtUY6qiZrOy0TI54BRt7i
t7eFnxY7fIXy9FqqIcXl/eZVEkjVTBTqPbn0ivaO+eTTEJdUcBKvSFFbNyhckHzX/0h89lnPyI6v
GUk/uwRkUR9/yfm+xTdAYX17NXmReSxgaz2wJg7VfajyzyjvQbJBPVaLvN6Ox12lQsB0o4SspuXk
t2Zr0J0257ZxbTdOKXTOcaaMMCoNRr16WRtj8pkOJ6kRsdlXeCeUgocVHgi91g4gti/0btp5SUeZ
ugzbwhzD1agBbwqU5gaxTCAff/bdWj/x/IvyU27Ju6G6JJC1V0HcA1L1ggUpfVC7zcv8QFZflk8U
qhcRCQMRfayg9Fui0EgyeAfiHPKwt9byfDR8aOsvh22N4I5tNTYdEVjSF9E+laNL5ONmqMrlQKos
e3iWUUWRfgCAhrPMz/CIUfBZQ1R/UByvet8QNyaS+uPF/XnKtq3sawwS32hq3+d8R3F61eBCvvBG
QtJTW5j/KlnkEyNQclLh0hVAMxZMT4WnEYcS5+HvxY/+9rd36rPb6jSzQfDWq0IfL0hns+2TVRHp
u7n9JwWCkJ7+NwfxgqRsKClTpzIlaT4CslLK2EUSnZmluluBurQeNRQbFapjUt8vei2104FgD3jF
UkO4yBZOkoAFMY2d0e1rmvpXgInaKoZod8hkxEqfPosOzLHHphx/E28DARXwGWgtoJwpH/XZO+rE
nalH6v54r6jKpTc/OW56aBTEETWvjDvciPpLR75Qw7Aiu3XE/O1LF/eDfnqzSSE2VFtezIEET11S
u5UJWCK/OP1qseOWegX3kHJr04aAMI5TJp8GDWqO+UgmuK6lf8UPImTM28/zxZy4oJEYdR/OAjPN
z/zhYSdiqkI3Y2Owla43QoNyB+uLGlsom/t3g4j8HMnqFY+/BUud3bvAziad29vCIQAEL39abOTF
YlZkuFYYq9X2FyEB3CVC5uILbIXSk4wvqzgZl1F7j+H1Bt4DJL86HZkaFOaGi6VAmkNLeUqXMPTW
JP+NoEGNdWVUyOCCjx5NW9zOAez5U4VSA7Xmp6MrNGg81k5bEi1bgOm7kA7TyNMP8d/9ipZyT7Gh
WQedmMNPwdAafAABJE+aKejdpgamLGdrXZOzoEfmJSQg/afLzu8bi44GtXp5aOxMnfiBNWslnGmA
n3oBNwQI8ToB3GnLY82fwua5uW7i4EwlEwLj9T7W4ni5tcl3VteJRYuqQ90HXp3Ml7EOa/CAVBC7
rhli+MMcgv25tZn+YKLIivgUOocGKYA/K0myjK0gtupgpn2Sgr9aVQzgYgmOhalvlVKVWkphVrG8
5pBWcUYpAqHR/IxiZfGMHwVJWkZUrLqCte6Oa4X7ULIwQtWSweo0eOZrz0BeyIhqPfIzgjrfEqCq
/JGuAKw4KcodchYjtsxYhocO6DdyVc9PKgpu2ZKmafK2oeXmM3N5t65A/q7BXxptuLi+dgocGoGn
KwextL/sRR7eXWqGV15AlMX2fhXF1byltyRXfa+9MizeH/0YMSr3cTpdJz40/uPM4tt0L4dd3gJk
pBm1Q6CXvJBSXKQW9dbFp6BCey/HVZrFDdfSghq/8npF/VIocx3JHvH0/yewiSK1Ds1yY41cqsu5
u4bo+e+Zuxbo60nWAOzTBK9ve8864WKtYD7QTwQv9hyjCM+qricqQyb5kR8Vy35v1tY+i9hdX9wT
EXQbEyFikk3TkfzFOktioTWVOK+Pk9LW0l8GDlrjxJXd+aHU2Ai5iBtsraNYXqGjWV7TSPD0uUuE
TZssmxA7qnQPEAMYVeiHPlpG+Ecb45GiAVa+WCzEu80d4wjAYEMR4kbWrBvgBPLX/a7eaixP2hmF
ydQiw33BEgNoL7R2ymeAPvLBL+k8J5Z8gmZvnpjBiOy64i9Ce3GLlys6QP3QGY8WiSiDTAX35pTE
50e7Qlh3oInzbieK/5YyfOjqoZ/dFPCr7M3jOV6sktb2vWUblPepdOMtzeii6+LWsDLLhG/GvjOc
U5bs2PrbdYKm3JwKUYvP19f+M6mgGN9zmbujUXxE5Dd6r7sr8dRyEsGXPCN3blwFHCgKHcrQNu6W
lKcO2tWvaAiOU4Q3l06ZVT9+ivjVBBgUQNe+4cgYYUphAYfQ2sefniv7XwB7R6DW5TGX7N+YBoP8
V3MrE741E95XXGRg1sxyn0e2m3mDgDvRl5Y+bzmxpBUhT0Cn7H2nPgZwymOWfUjN4btZ/Bj2yAw7
OFMtnFnw65mme3mR6wtGVPtJMJZMTHgJdhiZ8t8j3nPFcOBQ/3aJTXGM2IVHTT6/lfOJMmNCKDyN
bt1o2bFnn4amnEPkmFiKXkon5wDYAsQ2r8SboNWWy6D37EM2WQ3/Bpr3jq61gQdbMINdS2fnlm5/
X/cloZF/LNK098UJ1VXj6dfUGo1fvpMgId669bZizumGYk3qvFCBAaIjHM/3uz55r8s7myZRiesL
3nHzzBdp8L8HZKmUBwjTghWOiFwfC//6Vc+mCRSPctRmnRE0JVRk17m9VYZtghKMfjKIvAOj4Ynm
GOXiZ2wHvb2ilsnNgeKSMHDUge1vujqHSv+VdGNPBz2SfukT+5yJtA3QwVuLsmvKHd1Ep5KwPrbN
GiDJWXyQpdYBjXxdBRmgqnfodVq9I/KDVjI+YRTymH4XDItcwgmY8m8YVXifRlWD1CIwas4a5mHQ
erxFjWeFmVoJ3KFkQOLJQDzWTnYyZr8meNE3mDWNBAmUuq39e4JU04+idKr4nCkPRTQmneFwttfT
ZvIPYM85L5C1TiRUcRRx6SG4GDwJAbYZIYBVz1yiejKbSBHmv70QH8TW0CB0NBe8C6gw5xgj4pWg
J/a2vrKU4Ff5KKMuvok9wFQcnX9ljh5LKJdCHQdRL2AqcHlDYIR5MJPSVMzBjju++rois2iQqhKd
BCJUITa0K3aI1bataZeOHFNUV2ZZJAuDV8yJPmgt1zV+2fOjAhkMUze2ULUktXY1UGFDvcbnnqcE
z5486UUtJmOmT+Pj/NrSZzvxawwJUk4vo93q1P7M0IuJpXJIYPB1jAcPv86/uKbfxw/U0R+Sw/jW
MMHqZUXd6Ndf9O7FhaCyjpdNWsa77yd2A30jGPJl3JnPw2xaX++9VCIeqNoyc8N0G2p0vwqM+ZP7
H757JSKMak7icnpcSTu0mKZRxK3YQX+WazsfrDWmSqZaqWwWBZy/45KyGdImlO5A3gPrm7/vm/ec
5q24SkVFVD2ihMEfErY1uYbEzeDvhe+9RCmIiF07qyILkguzeXRV1YGnk5PqSOMDxw8v0fTjc7EB
/ofUjp+LPf0RpBvSU3frZS0XeznBnZ1/8IqwITLRCrSau3yAVWB8tocSsFxnX8ObNn9QPALd/bSa
lLgBi+xKvxKiHZZOL/YSRbiT7c3dTk+vqX8Ig/XzF6PBxaXa9zQxyGe9aagu4TM2wFkxKgPzg8+s
z+BRDwb2g4SJljKoh45xLLGzaxRGFXAApP8lWHkNR0St4+sc9KNP3AnbaxsTFCGLs+zZ9UmEfUkq
J/S9zPtU1ZLwgrEy1b6pPSsZ2oeB/f0bA1Jxz0MmWATouOsBPrImN//EiOI1CND4CAxHjD5+O4Rl
NLVGw4GIQOlAdLVnToxmNx0Fyx1NhXq0stIwcuLVvHuewvF13fh89go5Y4/ty19DAOA+G60W5iLg
skVkoVdFzypof7gDeZdChna2D4SWykTwNUsi7MdTsn6sfGtQPGewkjNxNhUNhxnCE3mCvDVV2oOe
bOFHbiwQFdCbsurPoeFi+4Bl/C9+D4PCC6XX4xEW22nU+8EeeOXM6Ox2CMrTHzntpgOuccTZp4Qe
EJQ2TUv/hBm6X+zrO8KHfJ4NYzia560hUr4dck88krsNQZM9uGMcZKvP6lTF811umlteIMEvuhBq
v2FkbeETifhkJZP30aUD+sWIrJraxVP8poVKtI9FThilox6XfmBDOWHoN2U8t8WkOQCGIZySKdS4
MJnptkwcU2w6n6sWsE0DQtfSZb7y3jsR0eEVpwUJYGxfoJElixrk4OlpD+1RExA2yOBA+ArusNwi
hQCzoAk4cDpZj5QsnLrol3JOfooGVcPPNV5X8qM6s2m4JcIHfGrnAZkVAGbLawtN9hGVmwOZHiX9
3oMLhLJY4e/xvqAXSvuynH6d+2q1CDR2qMdhDKmjmNRkutmMROw3EQcuTIPb03fYw/fqejtIqqr/
NU6LwIy57IC25GIVKPe/5FrjBOtfmbdbjmX3JBQfUAC5/o3nMQWLR0HV9cUmXF1boow+ZotVLHtm
8cuACLcIT1rCX4b5HHYaRvhrkHsu96zsfXH9lgE7k++X0Y4tECqEj3+Bzqm4ws78b8+pqVNnRg+l
FOZr2uF/0036LunowbxOfPMYdGTeihnZw27lqDIqum+8PQHiQU/q/gM5sAyGWO+kHQ+Rxm9kvoW0
KgHMPeayjtn6CLACoPFcHj/tdwGCvEwO8jcKtcRNJNCPo9MpvVip3YCa0iszBONxOsomMLjypfpV
7Lq4LHmASP+ul0G19AO/xHZde7WI/xGh3hSdw7UzfSOqME6UYvhjEzuw/iACl7RvWDTLJXExs6d+
FyunoGh9x4PRUlGnFctnaN9R+HMQj9/xd6LwhCwmWmzJwBxBpenxk6Xp72n8EmWZ07E1qDJAr0z5
jHkea3oXiDZTxfLbJRyKavrIRFQI2qfSPrSkRlUMxxSY0W5mrdpXbLMroDD2ejNEFclR3K+TfVQL
5mTSDQKfZBCtXSzcMH81ewYVIahGSbPz41Nmibc/ckfRRPGK/3X/kdzF06008q3pGLRDUKevUhH5
RIyQsaOyJ1bljnU6Yx0fcEpnE9sBpGps3DnyDKFyrLw1XZlLg/EwxhwGrZp9b7pA/07V2Pbh3S+Y
b+KP+5f5ZHDFUAivVoazEYjpNu+h+plEzCNZAZ3NKzNraDcY5OW4HPQ4nh99tR9abHR1mPB8wDzh
hn3ecLDaxoLxvCkY7Qu7/IZIrfQOlKVd/2iIJ++FIqJQQEDNn43qbZ+heBaBTvXYJP4qHrjkTmDd
qGiAbJbYUK6x0E2zH9hOwznFl2pCZepgIXW38qTbYX5Sn5Fy5mMJSDEUiqpzQqqT0hyPAhUUArDF
7pUvfk27/H8R8S840zLwAQGcLU1im11sfWwcBvEcLtDfqjGo6XFwU1Igq4crmxufxJvwmvj5bOar
qdW8N+qMoBFn5wURMZcKrFpzRs+YP1ez5drF3j6ccrlPPDbzGDiNBMrMj2qXYapanFDhKdP7kCxO
ihttRTRTlXHPTNTjpfC5Y6bKSTrv2MBW+hJSLfQ/Mmj5UV45h57eNqUKHvfZTbzVgJXbcLslaftK
nSWXrxhJvVmV3iDICOYhYiiFEOA9/pOIjzUNen/pDUD1blMyrCYnPvOHaVyvK/DZUAVecef3YVu2
k0vOOnNCWQxYT3kbQkNN5nDFv8JVytL11NeBc7qN+oamu/7btpgQJSHpXRcrUqD/tfPPu4Ahl0mu
sZd/F+AqVlIHh7wl8z26uhwp66B6hwA15kTa4rdpNWRUHfYEMqExtnKkYRysUhEULEC0TwrjPt7z
HgEScC5BgaDQxIzOxwRhJSdelWkcf0z6f82U/Jd3+T11cYNK6UEhTWUWJWGhdd04keuXaBdAwB4k
4znntk3jy2lrTsIEXUDkh1qfL9V0Xr60q98z+mz6RAvjCrIe4EoBtbyxc56DArMwM0s8A7Nw6H27
TFkkGg5hYYvozqqH+b0wvTBdDehK+KZNBWKQvE4pIrRh/Dv8Y5IQLvB6V5uIwtiBdtS+e83farf+
3vTyMTPeN46b42qt1wn1VkXjnGCdlXfcP5zSVHAcn3aYMkV7Uq6HSysRHevW4v1K3QFw8wbo8JIY
eqJ1ZlnDYkoNFZseJmX7Clhrpx4dtFuo4pLsvO6sYw1tjr5TdifJwLBoHLp5Cl8M20ZAaIEg2G3E
im5P6NVtUhFrmkXytL89QTm+3WqsBsKiVxweIgYUeSsdWS4JC4nDfRXbRrmjxrIVhlqnXSYy3FtX
u1s6IQDFy03ohHSiLbgQ4aT+zPIZFKc6SeMcq6p1XyWkDCYuY48XIRoCpuOQy4Gd2NaKXYzRhT5D
MtBVygKHNjGL/bT/BKAjXaCh/yPXDhDHObjMquXO9Dl/CW5zkK97lD3aHpDrsLbrknqHBbDFbK4+
KSBeQPxBaMQiqrC5t2jBBCBFrqB8KwBztWg0TUIxd/0M6BVM5VWnY7lXFIrMnK+IVTDbRy3t4ooQ
Qr/ZaSfDSnwtksUUQtDz9Iorza/Ce+OEUy2QjSD/utvnq5VQERMkhjfhu34N/nMNvStXufj807jq
BHkW+BJy6qQE3bNY96mzChtDF0aNcXXVw42CALNQ5Z6SjdWEYriIZvM2Rr7a8qAKJcGN9A9HPdyE
RtbAgzxO4zVpgaDXPjo9WGGHENdMCRhQoTapj1nF/ZK+yivwlHF6gQm2Pi2yJJZLshkASVsyVem8
TrAyAGW7Ely80zku/5w7+uXoJiCLn9Jr33dg/33q0kj+TGg2csVnr8izK3iRoABOrWSKE48sjhlk
t0qoL04rSJwLYdqZI6j99i4HpNX98N2akbbxfUsoS4YoB9A4Lem4loPKVk8To+/iIH1EbcRTj3Fw
h8obww9uvWoaaa2rpleAjheZxe4UD6pzQwLucs/eWYojD18vPX8oXRvs9f0z3TMfG2s02GwsEYOj
LdMjbqh3O1NI3vLKz8Tfw95IEaxx5JMbCIZwE7pdeI4EonERsO1+NQQ045st5qElZaLfxFhrS686
vt8AsmKoBFk97nxsig+Q6gy8d//QlatM0TalB/Z+23udtwqowDlodkkin+5Do0cIxh/6vErt+hM/
IZ0q69ow8LRmY0NX0PR3h4L+Ai4RXD55Kg3sCpCe/x8CeCT2QmcRldHNp/QPxlTJBUNdFwMsdhFa
8T8GERsUSKB2GmFxEdWjctiiMjfiAT6tiXSra7F8n7M84F0KWG1Tldoo6agytcue9mAP9SieX/Px
GbmslXMEcVw4dc4hucaoneoOTfbgj8e4XGAq3gIfJ4/wJ4hTYxiTZ4tzanfNm1Nb4/dy7oyzVLf0
DE3c6mF8HTpDYF4S2bS1vHXSqRkKj/4LRFo3uxie2L2UwIfdi8jp74+1vpC5jskjJxp9epjX7Ilo
SyaQ9IXISglexUqGb4B0Vcd3Gje5KiDOHaZdkS2WYFHJTDLd7q6HmMzzuJNeuZejBOilz0R8nAt/
6UwhwoLBAB8uoczNanjSZGSlxV30/UG/F5TQBJmKl2hD0SrpJbEP7lvRvJO1aIEsgvhgZr0eiFQO
/HEOaFphDm273+xed6XawZNKs5XhnSAb+ghE1p3afAXCDt67JMGM2gTADwdRJOMYLoQZ3re/if+k
RY2KyYHbQu9Lco2iGk0J/cpYms99AeQ2g6FLzmbbZb08STtTAO8YV7LGRTysSj585cggh6iwEmp7
sfQHzNkub1yP+ok5oFN9SYVonmwMQxfcdsMA6DKHVhVtyv1Yc+psoaJ/vzsriJYtd/nTDVmaw9sM
QqxVJv3eLmfPqPwfTWc0JoXlCcHfOAHdbOnKteu5V7mu72Fn6TrIX3C2HSy0MWUfcXbfA2gIcC7X
dF6Uupakc25w52sGaKs99XreuLov6j1wChTOSdg65idYmhwwdgbN4rVnlhESnbvVNWWArbxtJT9W
6y9pgXojDB4YsPS5s5U1iUT4/CFz5fBX1sPKVMntdn5KCMY6+xOH/M8OtMWo8Xp294wVUJ/0M553
8EKw0ITLRW3p8q53CigH82MemJ03AP2NZGLwYY7xfBsbm6mJhU3sV55SQI2JgyIHR3EIOtOHItPB
qkJZ1xSc+WrtspBS94LUT9p0fO9Sk5nentjiMLEkiJ1Kf2QKmACjvRcA01Y4Fh2DKjpwzBwrUFBY
uPtPfC97jIsPMgvBf5z6LFfsV8lYV2rucjD6I9UO2U7Qbp07fwrhyi33cyqKBN8VqWLz9FXCH8S3
eybZ6YoCMXXokaW5JyVz3qZt6SKqhMirx/xbnY06saNmZqMq4uKEdC6aXOR8R8ehGwhXGG57wzjX
8YLjKUGsjP4VvZ1wGUIlAAT6REhN+NLSbIXQEdyCDF025zS90Yi8DoBRD9kI+rVBhBIB4+urhpFO
u872qcO1I51IV3OslRvQLBduQKZRMBVp3v2EgBBPJ0Cai5O2S1y+wCc4r+L6bpsyjgIsnGNEqLTU
GoItvs2onzG9V4FcKmYJ/eYfnPl3gln+7TFX5m00skPc7A/+Ipcm7gXh3vd7Vgc11mTTVAzbaf/F
YW7rp8Zff4HGRJRHj0Xjc7OL0XUzaNI/BLu4DOgRLJgRcpceVU9OhtSNZ6eetRb+RY2yGuHUSoWH
Kd7LcJDr7gx9cxu492q/BAKAGgneCMJ+cydwPeJ6csOMWeY9JsLxdR9r+ZG+RcmDabqDMtohuaRX
ggviaaCNvdRce3ckhD1iiZyioOrT8FWpfumb/aRchPD7CxO9j4HM223qjuXJgn3VJkazwuma6kM4
PU/rthFaYrcRefGJOGeE4/BOJOzcPPCQ1DGltv8C3wMhKFLsUiUelxPhrDFPg/aqlIDNr5kD8S5P
j3ZZDeijn8DtqJj+M3p4rHisvFhivyFjM3hykkyPEjutWa+ARCidPPPL8Quk9oG66i14jy13pxR7
/K6f/kn9/zQUozsVzUI/I3jKBzr0L8rXF3dCjH5yA91heXY1LCIiXcIqLmJizdTeTtwKcEn71tkD
EJKmKtSI6Zhs+vyUm7ZsRzmXhj7ytLaluZQBk36d2BHD8E12N+Voz0HSZ4p/1wP8iYxrNYHO6ajm
Bw3p31zhaamrPBGHMxkOnpZclDRVT6GvcRQZa3WDPMOR2ma+jcSk9AE8n3c6ZVdCNiYkceOFVjAo
etO8NCNCWsGC/3qoxlP6z8BNOww2rYu7D1utQkOBUzH0QzX3cBsahiqoCqWwaSXVItnCliSpKLZw
La06ZKu3k8dF/zVQUMa/Y7qJb78MwhnpbTFXDePvPfwQ8kEZ5R6kwIgK+QwS8QgCWzyOfP2qdAUV
03RUJzvmzNYDdb4N1I7aCO9siRFaAesVaKReX65bW49S2x6ViyzKl3u9J59jfFU6ddY3Io9guW6Y
3Qpi7JFQhIecpjmqQvMYB93t1b+ELbl5ZJ5kgIGieJk5nrYqgarDQiE+eQKZydappqdIICeqtKKS
+dlm19Xd0S+A0SWUg0UTwijFGQYqfYz3AbwwbjSnbWQfAzcEFMgioeh12SN38M6BstUDfilz7rOm
ttl5B5kNVKsczpWXsefxLySJK53U84r9oAP4wz8S8Pl7h7sE9lSeybCgYzbY9hnrCd/7ehyzJhgQ
Wyps+a3ai3iteF0w4Ao8Jzvbqk2ohAedEeI3b2rJNDLUaxppWO0M+i9ypw6llQcbuMziJhFIpw4p
bGMsOq6kW6Y90cQQZmI1u0X8nDqtO6MHiR7CjEcUpUBDzx2nbb2dA7909KlOxeZhkn+3ryOwIu7u
gz8kXsaLvgRX4ZSmTb7moLit6Rwi+00AC7zolysWI+pqj1ZNjfsDCKSjd7qgBDl5TBfMbOMHo2oA
tJllTX+PitZs64MTLIyxulYTY5JlbVB7B8R4hdI7pUoEBB85w3uKWo4Y+m1GSbWjdIAED/nEXzZK
pMauLgtBFjoXJqEJWP2y2riHFiAJ8Gkm88hDcVY2dPUFAG0Z7GdoCRtDHc9oYzbh0EiQZQFxq+lT
YAbihvO3oNaNR8n+tMPLvZA0tBgpuLny9P4iU9dsjTJmu4RrpoXyBs07U4lf/YcNrbTwZZn4+8iq
OTKQUmQh2iqow4MXsgtVMmHvfO7UxHb7KU+HyrzdWpoTpvE6B7b/CPR71ozN4xHKGtQQfDTnWlqp
ANQtKtCsc8K5ajPyvDdfgfCb5vDIMaVk5chInAlqgMm1bvSSmEGUoZQHKMfvOht+7elhls/yPK5B
7FRB3T9rOHE5KCBQ+QQutcliNi6B9ZOPf9pjWQtQiOIFOPhSTpYD3USYVnjk7HiZ1kVS3AU414FD
3XE8cXEaI4O4KL7IOp/iM0qOfyvJqDcxpGzSZc2Q9PgotCzLkeiqEMgqOTk75Oc7/p/KTzlpG8yj
4TP032YlW7lnuYv1Mor2RqyX6Gf64n0TR4hZQ6tN220NIp0evYShSqwlUxlHXmNZSSJr+wMZ6mpA
jBz+Eu3cS/VyNSBlVhnZ0YJdxE+fBWDD4c1KVjYmaoVVngKAFLQ8PcYDXA315XJ9AP1lIzSmar3q
VbPz71PIwWZpBPiQGbu/tiuXtm1ZAWEplhhLnXsOGcXX4qrzZhA86qi1B0t6tTJFBSfSKAMoDF55
6QmRKDF8ZzV8pI2wHnzOQnt3GsTj6xJsG39ZgSRrFqb+9COlpQDiiFHgWti7P2H6xIjgz9BQcib9
Mje/Ni5lc7MfLpUSGUQhe8se2onZ7E5Kfd9fz+KTsZnM7hVyOKRc0Z+OV+qZygzkQ0oeLIhAvmOE
sSZqd4ZjkXO0b2QYtGLJC5US9sb1n1dmW4YvW71kPgnkrDSlQ8lucqel/B1PYPPEnQtvovy59EHX
TciYirgcs02Ila+mSdaoba9lc54Bo6mXNas4leKv2jMwV6oooWLq5aKjHOtPGuSClRBP8NVWAgKb
Rb776+9ju94UEhsdoSyZkSTik124GdfmCrpMRRESe++p4P7eUf/buDPIM00MtfX0+3ubqrP3Vhat
PzBZbXWCTSXic6UGUNBM6SW+slhS6i1PZ7Bjo0pecG9BMS/ulLJIbZazxOKDX3carWiJL+MbIpi4
BfgEfCR/Fl4G/lKlOS2N9do1lqO8ZlrBrEUg0jmoy2rF9lVh3wvRCi3sxJLvJ8KigFH6zrIzxZTg
couP31IyIhqxEG0y7W63x9ES8M7LLBQGXaBZahk4BhpXY73OhmHi3CXZ0AJwNbjmcAPZ683TMbeH
SHphUvrrAMwmnEbjM6nruIFMyTHubNnAtxf8g/5o5qPKrn1yyY8l4jcDhmzzQYYQ/H8n/YUusan/
O1IKBBQ/jiKjeLj4yRkzbnr2TDTlkm5He/YxLUk74nKOFzK8utGUCOJjt3/UyQTO1CazbRuG9hwT
2OhHhfusqcwtA0Epa5RnAjEbaJXbOC7VXattGriblfcF3LBeiBUQLH43zumt7olRvO6LboUlAn0s
LXsbuJOt94+Q67ED6kmv0Yup/pGjXRy7jhXEyVfJ2wsKdhoepLUyOz3gZYdISsQuP1fIbmPafTS7
02C9KXz33JIgTbJfMhQx6yY4RC6tQ8RuheRmp5XeMqKSs1FLD7JMDFRVbD4UgeJBbQ0qA5lIhZ9s
EKMUIBmnOTqILfrgOYtOfxSaldsOdI43EENOBkb06QhSe/IhgqO6UBhltLbsXOLzC3yc5gDHEHLJ
gqBt0BAw2BfQIezDEvXsRa5vUEeRwQ08rrdl7BJ0PQj0YJf2Ql52O9XnmI5+nNVZZrIxxsGdToev
rUDIStwInAKxAXszpryVxqlsXKX2aXvNrOmDkbjr/xO4JK4ymDLu+wgS2B7wM2oh+pkf3Y+wgCaT
bGnb4v316/F+opVdMXWjXfHnDdyTPs2JNWw10AvLWexkgxV5i4rS8H2+dxURzk3Sml16bRkUNnf+
zCWcox4TaxalViuAXrgaw/DWSdrPdZlAs1mrzcMSUVH0QAqFz88CgQhXg8wdG0Im+QXRfCHArX7H
TeQfe+vV6hQT0DgFJQ1kvIgfV9YpMRc9ruo+Zs9QJVMn3jyIAPIrPPvsVeFLCsPVB7FzPeSgIdEY
DHIUubzM6S0WcMydgNvn0PU3cbG2r2UUuO22lqEkJFRYd4rb5N3BMaa1I2Nq/recMZCVb1MeKVkO
xpen3gA+pzP7phZxdh7mC0Gb+KEu8TbjoMspCn797sGBlgz1nvKNvc2aBc9CvzcVqX6VcEr5Tf4v
naqealI07fE4ZPELlWT/Kv/33GWIN/Ip0QKqdXdXrdrGzyK2gqDZhBH+fZxNYB4DNAovaOImPCVg
nCWg4qQHxKfKX6cn4WUVbHKzzuCL27iQeC19M+AEj2pIo/oHy5JLsTQPNnCQR9wQifChGKSH/X5o
Vg7mzLvIkjkYkPZV96mr221zUjRw1fxuHH4w78KsA52R4yOFtrKJXyWiRpAFerqQQ65cYjD78ud9
thC52H31brnUfuefejH5h2AA6pAPY8gb49il4MRcjEdfDrexwbyDS3vKt6CPw0kwmcLP53KCpjrA
bbIIP8orfyd8HhrEyWH2DKUHB0bRvwDOplnDK8sRGMaL3LqEQaDi/Rex9zbHehwk788EqdtaejUO
wtIK7dawsi42mP0ZwFhMDFGL+/SNqlyi0G7rJKF9nKdWNfMQJ+Ua1pmsj78402HCcf+PG7DqgwbH
zDh/GvCrrcZ2SznQU6TniQ3xgHsIWOeP4pQJoOysFSBffJ/fKX/8rR+BIjPv5gZi0AeZytTSgmWV
DRkKQ53pMQb3h2hlJ6RPXyBUfRGJvtvwLqqtnCYMmbMchNs0H2OV0hVzFCw1SAK9e6JFEYEwIiuw
Q+zFi0fHQfv0J6Yz8YadkpPRjNrUNhNG2RisDV3vZb4eHeXAlti2leoy66TxbP/1s4V+5GywRyQ4
TrICFxEgZQ8VwN1HfKnZ54RZApsDJ72gDtRe6JVn3rpuYAa6R2x4ENa4srPczALq67PAevYFnIly
Kob8DyIPcUNlaw9QKRrCPqysXsTHTOYoPEKOf0f2bo7AUsyOzjdYb2GYy280C+W/mQNUP0IglHB6
DRoFLNC+ygO+e2t7LEH1FwqyFX6s2JkrB18cTL3a1GNM9tQKQOzzh6Xe6qS/M7cI6BTygs9tkhYH
Cv6GIsVKt/jq9fw40qiSkMRNKE0MDcwis807HbJKgsH/ZpKubENJv7uYnIO1QFdeN3v3o9dHF//U
AKIdRCgXbT61lHKf8FhyANnZFK0pcfMPtO8L3Hmq5QfrQkXlC9ITalcAl8YOx1Yg5cKWpqgUNyqH
J61QfKnMG0OIpc4xZ11ZeOpSjpyfnof3lHxh7PIU6P+exBHRCX/qMxgGuczJRF31AuH7ZuNNoKGi
YiKJkF0dYcvEHqoeFnnuvyrBD4GfPGtfGp+y9mMctn1fKh1lSH80dSQ5IDQrLZq0rLhexfVOcdDC
bPzopvSPOFbBa+BIh+49ScUzXhSh/qGYeF09TFRxMtHonzwW77xd/6PKz4n2AZmhr2pvU/0qbrGl
pDboKm5wouyv5vj4dq/FKmD3XnhwVYRGfuWs/yU7fB61UNBvzgJWDtoPklixFJNCkP4YW/61YY09
7b+5d1aaE63XR4+JpkPXQZmvfXOt1L9RpI3CejteehMCovQN2weYklQ3QSBdY7C3C24KM87DmggM
Bn8DH4PijYbHp7KYUI+JYRg7yfKd41FVzTTu9x7mKxVaQrhZQ3WMV5FBvD2YtmAigIXhO2G7yf+P
6YoENLlVRGHp7kSaX3d7/0GxB2mmvNUUqm6X6wVQ8ZS0yQFOXvASgJcB7WeKWsgI9lRk3RMlIYjC
74u6uQBdmaasB/g656TmtymjidwoVGpSMZ25CfS65YYZ6I3d85MoHzSgcQw4j4hvgnH5HeE+eFOl
hu9U+i1Vy+fQSPGC1JusKoG/PjfJvui8Wnu/p4BVOJVjIa342jnI5TOZL1mLTM6AbMFaJPhiiAOe
n79tXTxlRP/agItjFLCGvm+JWs1bKKOW+O8oFuByaG3f5L8zPakoIbT966RxQHd1LLIM18dA10si
Q94WFWj7n2TICLkmFjDst6EO0fCK1wP6YyCPhHZgid1P2dKQUao7cpI1epynnv9vi2bRCAijc3Rn
QnuGUUS/C1PLelmGskMxPcvoM1ScTKcHtGfmAaZJfduzBfZXcliuboKRUrSit3RAMi52dF9b875Y
RtoJhcPDqyeLzbDnYPC1valjt1hE0MonGGdIxz6C3AKK+cwkFq46RvvDhs6bRj94UmHf0xH6avW0
dWuNPzHkxg+5AqnjEuRQDpTzxouckJ0wIZ3sHRP1OXEbYd6J2P2fzNSfWLs6XAGxNcMKL9gp02JH
QRPeVxYyvvjTljp550p9mHlVYZZkpIHB0Y/kbZPyNnbUUozAjmmObVK7FSMsEr3O4zKLcDvmH1Re
8IXybE0oJJSpQGixgXzDIGxxt6mjaNtSRH33k7tBHiDg+39hSpPdn+o0BS/MdUVYhzEPHJnybs8G
RouASn1ED6beEITDzoafdqnP8K8/NGik0t7KMfb0Fbt0tX7FUtZJg7xbdR7Azk4AroqqDnR+hpiN
mIcGEvf77gJktiY/qZ9HMfP+ItomCk40DQNIlfeQpQrpP8txLrKxJimVIsePxlIfVr+vJ8N0fuso
SfcKA5hwxrQop1UOdfqMCRiK1pCK6SUMOj79Is/LkKOzJX+nJUes4lIIid7xzwzpJn5kmBE3k10P
azxCl5UNrF8XWH6CIu2Z/yTXw9rcU3vYhPQQayv0w4D9M8nM8TIvBFEefN0lBUsmUvO0JfXSX/oi
J/kYMJBFXkEtXhfJWMafigkkcBnpSH/RBT/WbCYPsvyiUNQ3oOuWLYCLilfulhd5BeK2dYkReSOK
WSpS35jtCn0Xj9Y/zfPu41sTlNxDOuTSBi1UkAHAusmPJ3pkvdaoxfmaFVDfkufFhMT46pZ5/zlH
aXT9MEwcBzlq/NUrnZhWo3RsCyfSUW76Y3ME9TDcU85c81HlhIYenun/8ebigfLqVTtoCSKZMqKy
P43U0eS5Ez7zO38YPuzplQA2i2ONjgj3bA3+ILK6T2P6YqfHn1cQOA2m348Jshy2xlKEjj+bvlAm
hx/RG0hbvXiSCbJfEyUYVFL7TNXpSJLWRIHP1czFHKTGLlTSrQcc9yCTH+nM8UmGjMLMiggwD7/l
nfRleWfu/mXi99Bwut3jB2fkd7NQeRjP7l5kMwGNMLsgavY6kGtibOPGTGsEn+u98BxoInyFD2b9
Ou1NT59q5UixItUE3xO7GbAGwVoCihEEaxi76fCFGwhJd0vhjovmc/NI59mLhZsebP66743WzTaU
+A5h4gqH6D1X0KQOKyojynIyyD6GenASfHUboRzRNCojoV+XlgK1NIvHsGorbL3XcdiliiHt6Ovc
kHjsaggq5+vxd9XYOj8emkA7/TIwJi7gfKTj4n6oTEnMjvucWKhJr5faoWGqJ+GER7GXa8mAnQe6
kmAjhjGKefaeu49o8OPP5i0em/d0OjvFc1tdmP7dUC6OOzJz/xE2TrCMXcG8uyXFKG9Fl5lY0Gst
KuxxIxJBkR8XPN5MiqLGLpBtOtzUEL2vivOq7GREKqbPiJYwChRnAtXyxjmjSDtYFc2Kc/aFK65E
1IuKZzntZAgPp8UtSd0H46r4c514IFOd9nE6hMuSujvvZkmDUIsthMJ4OUOfAkEIE1YyHVAgCixh
k3cQbSHTfcPkgPk5jj62bPmJDbyaMyYuFyqvlGVloM7BlCX/eCr1Yez3RYoMsjhH1IKggw8IGtcQ
xXxGnpAPHH9nkZ1aDNsgzZzW22hHgLOodxLihedCPaKWM8orNSQWvLM6ryTTTiKS7KEaicexvegs
ApzJpLZAtHr7ITohUQRKv1JMA8Bm5GiT5P9MGTfMBNMalSinEoiOMPGjVOAhi98qRFZrKaclQNnh
/9bvTN/Rbhe6Kw6EYh0vmP4Z5p7ioZA2wDKgfjo/C2n/ESP6qzkuk8E5k6MaEy+KU7Uc7DhUQ8ZE
HK7cNEuFFL4eOOdwj3rIM9ClR4/jaUWZKnnrunTvX16+8MMjF8Io4kc4d6fQEYNAsrJ0viPCxyeG
Xi6UWj7Ui9dF3GtEjWB6xrEZeGdNMH7s0qFaaGM2oLPu4FuGIjxMqQfIlmEDXJL2lVoZjbQoLvEl
qLVfMeB3ANGRrd67OIH8hGp2KG4ftBXoX3NkUWclIXiQEtDJHXWBRHVhWMpo27drZDHTj+4q30eA
Ny6ic4evMoarrY+iE+ug0+tqB9/5rvzaebDe/NRMsSMTS98dRS2QYIc4dH7UlwMHWHpPdksAlBjk
qf7X2iHd/qVOJ5Q/hbTJbR+LWMnUEN1OYUh5amoUcnf0LuAS3tzbP1y8gZm5qkDnhjSXJuPiFWC1
3u2BO6/h9ZUNXuuA4rkid0ESZLfnLuw2OwdLqgizCvzpRCMY1tFxJYjQC7zZTfZoUejVzOfx2O5U
JWbcdUJLUsckB0DvF+rIpJLqaybNZZAsazOvO/O1VaJDe0pmsSKIStYv1nqJEcSh3amzCCMtIDSr
+lQ05hzcwA3U6u4xEk7+UMfQ+sVUbFnTiUjsFBIOGqwr0IO284QC+5DpiZ6WIdidnz9OuKgA2dix
p/iGcg55B/yggu/rFNbx2gHkdwp1bguPnbOk6BtFAeO2uy48eFzGqVXwHZcKpustHZfn1qf4yKzc
svlNgOtQOiaNY1Paig+jGCTyNKsYjD6/h0JgUJzChs4GvsychnK2OhmDVHvcQu47p4xyC9VZkrVa
7sM5ZJ/Z5AySa1VhS/gMPM7AtDhSw+dnFNiCbhUA+io4y9yrhp4qtwXQrB1gzS3hHriC5rCfqvRE
68mmmVNFbj6UI92E22IzwsyOSz7QJDe6Z7lHkyVLSKfCwplqSU+3YhuEUPCXbHyP3UNnbxsuYu/M
jznMScsV39ZMfpAUV1jnDgrLPETyw/LZdr8lPkvupikxOVit6yeIMf+SV/tIFcsiWw5NVrPxJm0c
anXBdbXsPgJ4wwE4+BTNR5fET7fQ0hoVyWNiXcGlhKv7FajNTBhvS+Vgx3Dql8f+b36PvMKfMZNZ
Eh1MydlsBduacnx+mm1eFkuAAVDePUlHycbnPKl0uKQJXnH/o1dwQOs7zS+Fs98VyOLSE4RMhyCA
tpUaAz7LD+57aFc7DadgNvcR2ujReoUoytwIZyJKC0ItMjRb/qfQ5CxzYYG37doOiUW6CIPK6PEw
B0MQWNAIeQrIZF1Zjvd/2ETcLpKavP89kgTu+W61kfKiopFSfPW6Ojf0HInntEgBLZyaT5MJiTI9
PoH/Qt3f15tG2Hgzza9ea9e1KHAMvg3UHi6sLO4uy0nnC/cznYwAlr32cNmeehYfTiUGgztv2s/u
cPDca72NS1pZfG7/WgHxCoPjJtDg26gbmqMyGj5wb79iFS07exCsScWXH+To6oHh3nXAT+6F/GGk
ZRp/B7UTlCMECFqp0SJpBSQqlI8Ml/gwitq7vcLdqyANik6a4PsRU44uDwzuSYV5T3n8b0CazhtA
cjcXKjEiTW3QA323xosi+YeGhX+0FGOCP5XOWGjSggFrlrTTVXHyDi7aiuhu74AMGcpV6ALsKHWT
xvtrO6H7hi6V8h8aLbFSAeaidrYh4QRaYP6EKYXfgO+Gp0YjPFPbNGmUixWsVUxaW+Zt0uQ7Jypa
oFD9jn0LwlJiRBIUeOtzGrKaPyb2JQt2v1D38HGEL0DhsJGAxvBpemWld0YumGA3jAF3NuaukXzB
p+8YPHeD8sJJ5MVHEglPGXa2z5nXDDAPv+8SMIe9PhVNSRP5YJLXtaEDpIgLoDBmKjpD4mcopZU3
bs+alNbKR3V4JH6aKgrqlddwJEYanERDDjN/b006gu4ZlhqV0aDKLWZxRCG1IlGE5si+7Gk1zHQf
M+9bNwzutd+7QMngg5VL2XcU5rQykAk5Ut2Da4aA0f87BikkfD0xHY5GS73jMynJTluYsMiW0C1C
6MCfO/ReJiaKcpk029KsSYYJJ5G3myaouxUyIYLUYd2eMxNZzoSw2tSjoLfle1XakZMCU4E2kWSy
EIA6VwNXsS4mP86TRVOEuSisJrmYX3OKoX5cXY1I+rkAbvlgcXF6sgJ2KqXHDJ8KmbnBD18vXMpS
PhKRIz+KqPccRZr8S6KtwNQ/Sw8KMAvQ1q3dexE8Ua/uYYuN2LfcE5YLAm6wW+TOGJurPzyLUD3t
hLB6+lG9Imb4VlVtN7uFg16jHGZEJelv3k+GJNrhdm2i9VFTf27iaCilJIuO0Z0OlYhuIV/dV13x
qyAPjEAbnlSktOYCH47ssiwe7J8KU7KwaL1n1XamQe+tL9owxIzwy/DeH+Kv57dSE8AwbP5+7h9+
fHgK14iAjDKQQCcAwhQqXNN7KGeSp4st1sMZ3o+9C30d1Iq8BgHNaD6jXhPA6EaWb81KTj7Ptzo3
8/fcKygjqOcvGgo5wqlIVzojyI4fQGT6yPGwa1NCvGe45eE6K1jsyOqT61P4oX/DWnat2Bb6uc/F
E3pywZ2aEGmNiCuKJKYfkA+2O7J8shExA1QtOqpxG5ShGY1p72eJntoXwo+9yNdN1w1u8Muv/dj/
kEiLyT2tVOIr60RstRchMyFq2gbq8/sHdot1/gXayhDW1yXEuPG2Cx+hcvciba1ADsvbVbGgsBYV
52YC0dl5i/RfEYePIMS4KZtJ+VuhEj6ZLYAZxOGD2NFTadukcNE5sHQVxoyq6qAEfKXwlXlNPchb
VDhJSOELGTHl2YODGv3b1o30x4EpD6ND0N0MIqL1eUBjueN3ryoHVD9yIU+qNc23uE4FWHwvopsZ
8rI3LuQ+hD/YAYa8cjOB1z0WotjE8yq50xjsLnLCe+atA6oIPHzXIElr+qkYWJwPomBN6pjkTjic
KQCGf7p8vRupOxMj0LF4FCNgdVS/R0M8nzcNX9sjr8h27oXVfyesEmB29JstZP17ZNtgv9TuEm5x
ickpuXcpNnfs07+i/JqDlWfmFfNcNCusKqtrxFzX/WYmZG3s9VRMaHWspj0u6bf5QSnacqA2t13B
eShoizroOg0bK1NAGJ7gPNDyGKvxDkBLlyyKNWCHTYwLCWQHjlsRFhiMDzoDFqFiZon+JuC2xg4D
xg5NCL30ntCUVKI2w1VU0A9K3X2Ul8FhV4fosRV9jiJamr3N6eZMRCRnOzBlKHQ5ISDc3TdoGAiU
JlTt/A45rKi5mxG4JL31wgN9OuJUPQcwJFebAn/UXy9Fwb4nguFRLyBSExmIK4h+V8eiqHZj9XeW
SDtCSQYvVXRZ4xqXe62WQ8FqKZcaiE4KArY5G21PZFUGO8h5YAn5+avnT2oJxT2EBYmKr5ThipOH
TIJ+UEuClWh4x1omLc+dDDtSKENzkZbl+LYPi0LHIgcAnoBw652Yql99mTPxY8DW/dmziZQJmO8o
TJl3QAnUYAA4kOOv2zMJNIUvLemdi2WMtynhG/NOHUvUWlAh6G9s1PlDWwDIvVoN+rTcfNX4+SO0
rfO8zzAf3vhgIS1rxB/Em5TK+NRrEC1P7x1lt3yrZgCp/P3lyr2eZmq8c/m35eQ1OC+WE5bwZ53E
8wBM83NxS0RvC9QBftY5t1JbnbvWVqs4ksz63lhxJmmohnmCCA1XHeIMKPghZdjlMceTrMooIAPT
CmwAjMEfJ1+jd11oJhw+YHdgH7Tfe2IF4M/hzFxyCZlqN9YkzxT/86jF0z6vwb7RdhR63AqNjb31
eK3UZ6HJkyyr7nnQH0OOGFTJU6xiH56gYX0VRmr8wKz5eiZJqX3SR5+sokgM9W41G3WfUVA+PBqm
C3AGEYadwX2y+/JY6mSq1qGxpokmIz+Ehg4P210S6+1BwGWYGD5QfrcsW3r2glrogCIWkCSOeTWm
ZyezdyCMidxmYfWiRf5E4rL53xtftWKvMatjGuupMwsYS93nLexG20+vwWjIntRWXLI0VxPrOgi2
WrZqOeGHcP1jRqe4SnCuA45Y4xrPXR+c8A1kSSxiFBMS0GhVOGyPisOrx6KiOJYDlHTjKgHYcl69
fiPspZsqCgQzwdaqOdK/B6RcxWawgM4c12SOlYKXyOZw+1sI/fOTy92PzKl/EA9/t13MeL+MPJ8q
fkaWWy34zPjH/qgbFK6k+2TURrGoa3e+NrzTUOvo/EIDjPdPPsrC0IevdRqFLUNbZEVRrjNLClEM
Yzs7vzqHWbsu90rH9X7BgolDpEyU/APmp1WJau/m0GN7IEvVzLUrVGuUuZKqHhLzSSXlecMU9W3s
mRB1bzONiHXwCVxK84VBtzn/F5PStv/70yIji4NUih9UT7IjyxW8AOwJ5CL/UnMORuCJQFLKXLrj
tibXVDwr/stUqByiJAxKhNW62tw1viN73bKTSAOnD8P6LykVzFMzk3nq1Eg+YRNWLgqoMX7iGgnu
lIC20vwFEOnSnkMegd4NkTDq6kjHPuQ4r+YmS39Q7110cbBYDAKN9Tiv9OBDxa+TV9RSxaVKFWK3
CIjjsbo7EchbtY+OV39eSjZsw6NWoCUvqHsnO9RHPLfJ1iPcx2hSQlzG1Wj9xXnQGYDrdqbPMwSw
yfrEzAJhtdLj1B3NJqRRJu4KglMWwOShonqiWeN0PW/rylF7tcySTUoTSBnWdIroe9DtLbe2O9fj
Nrm6tV4/Rxl/0gkxjXkNg8Q6jrtdvzfU1aU6lxTmidiqfrlrfLDS0AzLq+CSXSMh99Dg0YHdztk5
gp6bmRk2hmDSNOmPpRmdH5y3g2pBVWA8fXj+nBspBj2hSiQOIj5bZJk49eMVhjT+G3uhC90YkcFm
sj2dEF6xT1vLTNTZa3IocPRh8ufQ2IMez6eqlnsMBpfYqBrRqJUle4jqnB40uN86XK5QywN7kwi5
R+oE0iqFFnE32REotVLE6uL25TjU03GPGudf2bCKovNG6VHWw32K4iNgxO+c8ocuvV1Cw+w7j8TF
ey49+b9LU49TMxfeoJ7FwpMjB1A2fPmsuDJ5Tw8aC/bVLXj/gyItTvRs5hvoUqCdZfCgNSiDe+HN
Uu3WW7BQZIyBjbZNJUhzKE9dpWp8Uf1zAWpw0gGKZMMmxhkzXClWbLNBOEpEs9pJPSWwtx7YFBR2
K4tv14ka/J+DdL8z0QFjXDPvfHxd7r0vOJ9ZBtWySD8vitWDd004iuCdXXcg5rUDkHdwuSF8Ir5m
OkwXIcmk/AiwF2lwX8w/0jC+mvT5ine4RGnMOYX894A4xlEjEZ0KG/TcD7bLPRY4Z+T96eNDk63h
vd2h9vfoPsRKdBKtnD60y3qXgXv16jcgGoIArP1vYrJddNZ04bV16rI93G/tKkyN2YurSpclEBGo
wXDkOwP+jLjolusLBZgh/b+G/fBtZqLlN1Qd0bgu4BZV7ALlD0ZKf4XuuKSwh+lNsZdoDZ3wL1T2
WDMYJOyMvhLGLy73Y0uSfs+xhIh7toOCOzCQbXU5Bmke8n3zqbQd5z/lSpW/rXyKfMmOmIyyohri
Qc6JLxllBtK4TcAy0cShmKl9dTVkyoOn1yEpyluQYnPrXMuyWM93dHPTqRxZQbPdEO+AJb12wqxL
ZerzFeSdZW/wNk2PNmwtvYnCCF/ARjAPYyzn2Ckre3l8F020Cpbfn4GnL/yObXJjN/kWGJigHtda
Itv71GoaCPKF+7pSjr10zQXtoFCwOXR1IUaa50B5EaBRjLD2p0rJWc9kdfcmFjzVZGxXe4pdZN/K
YJJhhmZj77OVunhcVl9rojY4mM/Ye4bP//1UJ9VMk66A0j2sXqaLhFdbcRapNcspH3v0SvshO8po
JNHeG1NqPXbnM2TeRzF5f2eh6ilt1sFWzC7xikdEby38lRlkK3IClNVJVSKB4Lpwb4XgEMJJLsl6
nKsmL/jr3EPpY8x/7Ba4CsvnCdn8BwmYigBYGErqXgheAxxDuw4UTABKEuUKMx7zejkPmSUUVL64
Idy7xsYwvRUYJ3Qdcjg9n5lAoxYijpWNseY/m1FQTx2T+ucJdR7Wv/RpT8CrW7JjkZh9mF+ipoAp
zTHGvcGPIu2BeM3uGdvD+9NzK7CvumREfmeJdOGXvKsO7/1jTb2JvwPmARU7ec4ucSUua0Ru2DvV
FXgVAgBvAHY5N8vgLjjbjHzwcSj10hRtvoWPxkO0uriAnJjXso5Cdml1sAC8SZLl08jr18cByp9p
Xt1uRDk8Yh+n2os19KOXH/M4rQy7q3VykQ3YFZxRCXjSOx6QxCOXsFSpg+CGtEcHgIZ/kTSsfkI/
DMbp1hAM6aQxKhT9TIWs8Fv96WpkX2+AlKgP8S1IJdLOI+B1nKaizozD+sAr5vGe4hRFOZap2BAO
u9NOaMIa120raPcXaVJOsqqLXNROZhZrq5rHHaAY2TUiUu7MGRLXLJQr+m2iIYcEoVGlsK9dekiC
WdQj01xs5ywV6mqszhUdQaXQQBGq6VuSDROAWlBl7OCCeI5CNPVL672u//+xTa2fiy1ZWEAlTiKn
eAElm1Zt2yCJIASdvOtZCNyBNA0b5TRZUzUsG1a3ikLA+FK3LevZPsWbcbooaD0XJAO5TZTnXXi1
pS51ldJTF8xsfx/GPk+ILq8zT7pC6bBKZALTIZ/3h9My29NXrp5SC3f2kA0MP3vo5JS8Wi2FVWQX
0Fo5cmuwg1ppnRxL5DE6t0RsZgEU+jxk+v8WlXsoZ6yERUank2qJuvAX9e48pslH+nCQihLpzxvk
JlMOZLufW8477F4vo79fUf5ZFK86tnLhz9lhii6XolDeR2GUo1+mRR5TEUpphJstYzo51cLbeRIQ
ZQ6k+ki1yaO7MfXi1Yq2rraU7UwIaNPH8ewvoUGcCdI7s4uDoOnYT8R5nufE/wXBRqedvEol0fiU
A+5StqhJQPOthvZUsDLtHZj39YKD4ESFZp+2ecmpQkiNa1AKfCJlcXleVMgmYdJu8nMHF+sMxEh+
eGyGbTxiHYqrKK1QWrqDRrAdwsyWQs58ThWse88J5vDA9dDZ3GZ6eJvXdTDH3jPU4c77lyt/GAQN
In5IVAJPAJaLWDRed89cS8Q5PawY/eGHogLDTx1PAPDpaJwCQtCwRNvUAwZcvJ9vGZpm+TmwdpCA
8Duh1dOx8sgDNAz4++48sRVJTofuU8IeAc8zb4GnzWGIsRv1bjkxVjRd4yD24YWXlWTmy4IrwhO9
XSDCzMeaBWwO55NDVjYJ9pKvXv4ZBILBP+fmFybY394PydWcfRQPA9ib/OhC+As6gkfbyfak/eKK
3jPZr1WrLQIutDLsv1GrIV4CfQ9xP7CkGVe/LiKsYrjeZvNUbb/stHSZMnbl5KtHcBekAQgaI+G/
PZnJFl12cxx29KXhp+2IyY3EvJbDQy3Jes7sKMUNY+hnZbMkJceTtXH40NZZdQs5iRItkkKOQVj5
PTLWCtx/XSoQcMbOl3+e23XgFhZcby2rdQTmW5TDQj8yj68jND6oVI++U/kokySwjc3vFqUc6wW1
3fbf2CspAsmxV6UTPsDvzf6vMsKJvV200tmrqqodIpQP/aJk7xJ8ERWUda09mUPLZu5x/qirzeZ2
QS1N1T1nyTcX5Htikj7/iekEwlU0y6VQWNbuS8FAh5GXhP67SY9QGi3RJ0orl3vVrKny+GqpBO1q
u8iKboTP+hyNgwi/4V6HqnwuGju/juPV9uiswmUELtomkQuOeYJI6IivjTsBgZbpo5gTpQBidSsU
h6Jn99eVblQ6RppDOjFaODYm8kBWipYHaDOyBn41R/6iZzlZqjdKyp7VNaGixKAzzMH5aryXpTpD
bfCKCdnWZ+GHQPE8DxlhA47cUrwbphFfI2++m+Wif97mSPGARn325nX4nor2G0NN4oosXCTUcoet
94qEJQrcGosIvMDRWY3tFcYyKSyVq8k4epfBk+cfI/C3TTFQ/hfh9PlyNAoBVF/GW022mMOZO6mt
ZMQoN+bVYzDplVSxMhFC5DVLtX6KiHC+V1aP4ZYskx+DLl3HX6MzRhxohN+dyXiOryasOjxeYP4T
EYMZ+xyuaaaWZvkwKGC+0DVCE1x9mjGBXid/cVlMXQfQdWifKyuHYlt1BsfruYzESGPUPwuTxuVh
D7ZMwoe7pOxZ8JF6tcSTuP2EeSaLBhA94EXG38VWmFOV78Ci0W3sLozk1EnpOd2irrxfRryotg7C
iDfVIonIeQFC12/+fvhd0gs1yj8/4MQJmbpWEZJzeJkT+K2CvsrbeAiFbpSRrCzBRgOAs+8QoAgU
uNLcU/ssovJClVTf9pXaBokwecT10g3qJLVo24cBpP/3OGEdKo9P1pytSG4REVX0cCaC3syFZ6xK
EITNRl/1Unlww3kbdwDy3Ro0GksEC0Oif88yhtX143O4HVm5jaYQptWvGCx9TagxicvGyx/ugMae
rcgHNN43Xykss0XKO4n2JtTRr5/4srWZiXSzCGE/oNxJd3WuXCYSo8yBfRMeMQlasCoIkM5KPY0o
6cVpbH+THcIIToKiAkqchFz3KIa9wgygHl1PhxFku/wEuA29ESBbUAwyx5Az6Lu7vENrHFKlx5Uf
HopOQMJBplIoIRsfwxJu0MmjDlPl8g+z8Egy4sngM2sScobPuLDtUB4iwRRBCDy0ODUKQ/v0RVLt
9eKQYMylRQOsKYbQEMkSqFW46w0CQvNIR8GyUNVN6L5D+8nCqwKEMqiINfx0E6srP8qYs36tuvbv
9B4L9ZgwfgQLExQ+JhsOUH3ZD1ElDUczsuMj3mrz5D7sNboogc0Enp18kF0bGTKyKij3UOw9eUnh
dYcyIbE+Yg3XvgL3RbHSChRila+Om0jPj/B0yTfwZlBhR23zh3Mjuq5P0XH5bIjzDlH3g77a9ljs
1s2PWjQCvjaG7S3hXeE7Pto3BopjJjvaLcII0S3A7KsWpc35O/V8wcjDpCQt1F1+uOuvJ9glc263
4ueI/qNJnbal0CvbBq+11gNQ1pfz53uxWg57wSb2fKfJgGUId3AWrHTXfhcbCKoqYtSYLft7OhRM
FDj6bJxf7WyOdPY2OKqThJIAHczFrKGiiIsS4UdiJUz3obt6F1bNwAz0WN4u4HBYtS7eHPcP5dcf
5D9uChbAE0s17+5UqmP+99nmIUBKIEdCAnxarxFY3jvR1lJUlya/To8XgGx4Qm31C+KeRUVRhIto
r3qiaJYvt1nh0AxHWATbrnYQLydYqZ7KfaNY14YbPRnRsortSIPj7Hm7+QG+r/RA8ShPm+sbB+dR
EJk4zueqfkOtU9CayDcI06iP2hljCyjHrdxOPOfRlxilzmnbQNIsBD3/bvO2hvY/okVa6LNCQq0f
gyKmKvNM0B51gh/UCqZipSm8hMzkbwQsGqzmmpxEapYmaHXVUoOod5I2lKIhORQIohBYVM4X9y5z
vk3hrLhI2HlpVHpuXmH69EgLoHK/CehoJ6Q3fb6pEK5glE52iRRzyVlA2bS9ocsXmO515g4RsbZ7
gPy2YOc7IvAnKvr8MUEhserTy5JyrtqKfuQnG4++nX7r+XlrpyRKjjR+tLirU4bYHh+W2yNOtOHc
XsY88SrBKvEbu3LJK42yJHs0rmwNdd9CmJE7b1xTof7bG6nNYsNV6jD830LUFkg9WFFG6AOwOxn/
zmiG4iFRojD4Higa7l4q2hAqVjQsotzf3IRJZU0RgC3UmXy0jA7QPmdFBkGhRB4WHQDDoQN9L9y/
C1B5rgULKsRJXQMktR5IzHiKd1YqR6WIMLFXKVaPyqt7OdtJnd+DN++/CJtRFmGL6uqkfC0IrmPP
XGUAiXtvgBQWns95lP9atKVwgcwg6RkCL6AFnYu/CVP/hd/hwoCEkGaiX2Cs6PFZsq/d4CW7M0tS
vjtdsspdko7IYYGIc64R7k/h3KSV0WYqGtMEx+7rFORlHxIEgUpxgUdNV+Av3QrSEG3cNeMJZcLg
/sZddqVUlRGR37kZoIJoufLr7XAoI1u1JfBld4dnMXUXGjxf1ulaPXeGEBO+NHg5G5NGT9QGjn2/
vWHdA+Ok8o4o87GDoexiiWVN/X0sCJyFZj48MOTxwvIgrzCkLHn+st1UDZ4pYxPvY/XcGQKwt4Ud
czGToSR3t9UWCfDnbG2EHAfKe8rik253HjHp5V6GoOCWhYR24ve1k7uKzNW2tJFas4q3RhJXfWzI
CYOek7AsrSBeRga/dVjmHhUagS63TcxqMPb66Navr1ckiuWLy6P7erb2hNIzERmRCxl7K1kR5pF5
XeABtwsofrRTnC0Lv+ieSp773x/vpLZ9+ObQNPqg9FgPGj0mJlwfUJJ+h9kaPa1lwjdanoxoh4gF
DB1fvqtZdIi+bbStl7FxmTsW03aXGa5i+wzw70ALamEtfC2qisVDK1sBmzexFfUkBU6VOdIVWIje
FMQNWKq66ZBzGyICcQOWlUEExBTbA0+nk3rZsKJLaHGnwzU6dg+4NXC8qQJwdO048LAdpZdMQ+Og
eKnnWOP/IUEZC92PAwRdQeAPM7UrRMk0juSGu3YmRG1GDNW/w+DXAdzn1mHaavkjwmkssAcByblC
QMANxquVyZB39E2m5tGf84aff2Dkgf2rYsGgv8Bw4AF7ptVGlSt//wLzwmescntv/+xsmUYfvSOW
o1Ot2mpm3XWopt5Lr3qqz+1OVWsDawd/QP8YUyz8Vgfnilkr6aQfbuKcPAA6HTIIiycCsnATMPzT
TDdL5crkAdLxaE5r5cj+b7QFqI5CCKUvcCkg7jollAfSkVElQGn8BK2IfaOZQ9Dpis+597V1iM4P
MmL0zsO3pYku5xU1IxThNHITZn89nYT6whl+mxp/VaRrVaOZr8W7qIIucvGuasqlLP7ILyqKTDd4
EY6MP0to3MAPB8Wo9Z0h1AzFpDLXHrJ4GL8yN0ZRl57dWtz3fxU2i3/p389oCT2rL+qieOfFUGH4
IL+kDrHcJ9TRyPRR5R42YqVxxXNfuaKs4pmgFrhWwwHZfekpZ5PmvksQWxn9uCvxQl3xZ/wHjkBP
DJXuxHSxbWnQcKIKi6L0hz8u9g6XM2S+Py5c3m0CYvB7V9cj1T/EYGxp/YJ3gPGmuyBnidZqbBbA
KrYqcukFbW+JOMS32wtOI8+Snj63ijWAt4n0X+sKGjtfrjTa3bxrfyjGbCQP3HqQAeLyrd107kj3
WY5r1gbNIJU5H8ML5GJhTcLW0sE3WlmUSA58MHnTKrPlu+u/s6NQa8K0mQp4wkTT+DkQF7mwRDVm
95dcpfFJFkPNM++1tLms2n90jFDowWlxKOK/vjqyWF3erod+uBpKjIYWicbiTanPQi/Cu7WHdcqu
Yg0b92Pt9VbdGuPuasW6/48868DxsDn1HPfKvrlbSDNFaZ61SGmN+PcQuhZO801wUNRnyPSc1nw8
U8oPOgm9ZSjHjaNpF+aQGMw7eSzCAov6dZcB86JBDflKzbSBFS7P95vmonZuclQl2oJLmqwzRh9F
gDJ1497MYt3IZYVCyQ7zIMPIL584HZctsorXB2+1csZ3nEhEAmLNahgIw5BOzjE4V+yTZp1n2R/J
cNohIBjG4OoqWEsyOrEqsnifSe+QtDSCNkeZa+kdCrGjrMihTemvpS4nbAurq4XnQ2kgfPMij/Wx
WUwLjH75jYWiLir4RgzoQVujjJrB2DaUhlp0GdWJO4ahHDy3ZvPabCVw8H6ViAM9XbwFXlNh5ZEM
t4AmHX/Js57vYgqoBkdBPg19Z9kPfGyOvDFxw6oE1RJjS3Sh+Knkl71OgBI12lGsQs3SwcOTUjRn
3o8Qvfot9xhtmT881H6kjqVcp4Q/wtVOGkc+q//4RUgsmfvgVQ0AKSZ61PWi+WtoEcDFdcWoGxIE
/qnb0bOyI4Gqk8x8cQY8pS5ajphQc6FlJx37DmfELPlBO9Mf0m6jqveZn3MtgVo8VZc0h2G1XX/o
x/Pv+PplbtxoXYgFuuL7XeVJctCwneuFbrGtDU8FtxenNCC2da8n0IvUcHCbbG/btZDAaoCeG/Ab
fUo7kM6aKXx4ITeJSM1pBRrGPAfuYqPYTjgb4KfRXvYzDJyn6galU6/qDzdM6DvHCxrphmM3r7SI
2/aDTMS19YwXe/zYkxOzhInp54lSJgrbckBPyyZjuGM3sTWXf+oyFjO5FMYRq/h1GTRPdok9h2To
OfyS6MaKnUjjYpjfNK4wN/378C2nLafuYqPa+LLCYoOAvKcP0KMi1ASxEsnt09eTbcb8RX3JZw58
/pfPHsV9Zo8zEmJcSntWlD308rX8hSRlt3S5E2A12R9bMM2dwxn15QCe2ileNuoWN6VX85UxC+P/
LNNaWiQ0AiVFAOitJGQhyaM9lnYGqgxEDceQr3QX/9UjkyXebksnNOwMV/YYP/fXWNOP7JFoDqqT
4nSoQIdzSxyYvp7KpqKYUH4Qe3xEGR22JnJe+F0Wd77zD+69c9fNKIYDHdD5twB81FzH4RyUqPR3
p/E4jHmJ+JrrfJQSysVgiodOrHkMYoqGjsB/A4htklqu9EMSlScOcpO79YUQlWuE6V3LHBYN9Es6
dFOc8blNNYK8YcClL80oqM6/apx30+J+nDEdkdcLkDkC81L+RCqnAplUpQjJ44o2WFA5rVRpwNty
kVyuMSVMNpgFHy2hCpbxBBUBXbgxAa2BQBErg2lVuLRXJGYU4/CWonf+QPX3k4ugRMv2zfOJWulJ
GCKwrcPU8SzdhJZW4XQP7UyrKY6xmDKeS7yreCu1sAoohvVtIGJDEUreSX7tqA/8eScoxdN8wu3v
KmeNaIRJ84SQy0icbc4//GKpy8/47tLcpFh1fgbjf/PjUKcRcA52/buuGZAt5sk7HK1CWWOPLgXs
x861Ac+G8hU518rwfeyIhlEonEg7q+792GngfhI0e+WoZ0D6zDJFJr4m4NRDfRavl+p74+q+U/WJ
aaPOWS7Ly2IcURH/kPeK8qvZVB/ZLiigs/wenDFbstfAs1CaTSJleq23Z+4ZTki5VgSayWOgGW+y
RHwCsgQ2rTeT0r3BNk/Ljsj69t2qk70o9JRiNc+QmButOFQ4ZE5kfkcULrItDm5ZASXhFRNvKjhj
802Dpph1198h5FSUJVNH6G6o6SfNjDOEb+1XWv1TD/qCpb6r2j/VjRvGNQ7xnmF/z8EokCnm4a5G
43ml9ydrh+qCxujv6HWyZSnbNEkmJcAEm9FzqyA+Owak0rIVs3xa6O60/fq7Ml9zya3uvS925mUR
c/qWd9BptfjKMVJbohnSEav2oBdR7kKbxDPmJWP0uYtQ2Bel0r4+99fJ44+7W1IlYdiynEmiK+iH
3f0K3g5nkQXkWu7pIeRw0IrqIyLW5VWLk2jRieJLx7L+5LOhnh1VEpziKfqgM05w7psXsDR+bIjI
2WRf875vqAtTKAeS3HDqX9sVmT3CDyYjqdM/HsOpgZVxeJ0OtDjp5L/uOaapxupJfPur8EeV3TEw
a4jQCLHpCG1t18DUB8AUy2VBcW9G2GtbPdt3lSBGVroLoVnP1qNRdxJOCAQ1c7OHxz9nECjO2ZHg
en5FN2xm/ct0iMeMSqQwWIKHgoc/8pCTtz7c7jVDNiVp+kB8nkivdHydMk4EqrB04nqerbIj+bkw
DpL10fXBgDVdrids7trGUzUyQEb1edSxvpFLN/Z+tm9VHeoUl6KUdwZbjRP2yf6XHvSanElqtRNw
/o3UpHjoMkOz9YJF4m+07zcgKE+FC+AtmTpFkBC2kjYfS0vsTeAb8gK9hiqNiEjfH3EdKdSF4kEe
glmYD3V3eZh8GHdw+zA2YR3LBJr1unFXQnIkj/pIl7W49moFLrC2L8jh/hM8dfvFkbG1v+wQi108
I5NFX1ISSL1xoHAdT+jIPs84M0zewhJ12Xf75me7A6LdRYzU4/YFyO5ISHSVgW/akVfSrPxa439O
BysVvqbIY9WHL12GHcg0Y1MqVG302Mj2iPTQN1jz54G/TTSXMoHkfwV7yaVPDcV3VLs8D9XsByRv
pXYD3Ng6ujKSHgoRC8RtFQA6sd4GoK6xlxVFVHFXjAa2HcmS+3ymdR2iZI5y9aGmMpM7QQmig8w8
w3O1DwvKH6ylhQtgX9yYoGnD3WqAr39sCzm124TQOy5bxVwFEdUk3aYiti3piDv29fSCRoE7SHqE
QTKso0lTSR2625qiqeftSNl3L5IgES9gWlFEDn1GFhL7r8dQ5HPEThjm2J4wFl6k7o/QT32wWOZf
UKeNW7z1hIiFOS3wOPCnBEEURbctP0XzFvr4bVuHcT1RMGB8BeaHQ8m2lN4r35THtu8lMI9BEY2b
bHQAyv1x24cVuWKCfJveNBTecKr3ncB2cV6/q1xp46KhaHiAuH0H5l/tQlsE/Mf1MJpVRH8vCnXR
gjhuanXyc6flkKigLk8WGlTbg5eNxc4ylFB4BFSvtNBiQ0iMh0c3YmsV2IS+cHqd9BUe0J24/j/s
tfX/W/jEUcFV/bBVBkam5IhD3Fuz6CXXsVoZp/HpPWYXZ2/yNLCcSA3CQNPX8FX0CihyUEXf/NQL
Xijo8kU/IUNN75zQcbw1gBQDU7ImDFeH0etYOGn9yXEEKhZFibZD7OkZLcQWDcXrVX/jCY4w0/bi
dU2bb8PvAg0w0aioFAlwHFBA/IG5V8CHOxJsEiT5GXEHrcRzphfhQouX8iLjdAqXIczrOzsvJLEQ
Q5dvv43a05u/1c0wp3mS7flUbojRswiY99mNOeblDrcyxy4/FIkrY6ApslxX0Wc6dTRcox+4OTbf
DnImug6+Egmm2yssY4SxrzK6wrCYHUfPneY5aG8PUymJ3+cknLNn7nMOCRl9+pEFwDtlmOTYsffO
wFvm8rIak0jIvlbDw7f2GV8Cxlf8hSEyqejG/BCYtQ/n2viJTw2x8P0nrNUBFSgDkG5/fBIU5Kj/
EwALbKZMSse9Lm2w6iEXiQJ/jgzZl+yWZABmarQE/UvIPT9XLdrjFjmG3fRXBY4TJ7VAlQcGp+zv
wUIv+F5BqCDDk9dJcxwOlzXox6QEhLrmaD09+LUtyIABZEvjnZSzON5p1TNc3hpCGMIWile0uYH3
BZ3JAFfsax2kcxZC9tkVINnE/zI9h3U2cPqE70daZEf/Y2mnxZxOhS+i/nDVxyxkdwLTe9rtHdCO
ftAGAtvgg7YBm7BWCCyRYA8r8iSV/3fBtWwET/zj7tyIOar0Lomg0/Uc6kLSWOuIoI3p/NAhYC50
AY/TYdJSXSvEvbjJl07JSBqmHWDeV84kXqPhox9wCLvlNv061Otdmv/Ggct8Olc1w/jonR94h9jE
VkQSkARPJPEr2WZMxhXZdEwfTsaBFwqF4PL6i35rUbCsav+5qWrU9Q23/QTuKL4FHfUVZFX2PLeJ
gqyU7JlDkK23kqD0r4L32UR975I918Dzf3X+5XEb0mcfhUbGo0/HmWgjqUXYbz4AXLiEjyZLrc7v
Cxr0XTSKNpCu1z+RFMgCilk4a6iQ54M3gmuX7j37N90LstpifNe92OFcxouOOzAB0It2zdID8U9j
EN1gxKwLtywfRi6SMH0wu5XEuzhq1dejW3QdLr94hK5+iZKltB+zLavRLY6BxfXwhaNvOBpJAAKF
qiQWH6JsYmV3fgNLaSs4x62G1KJzXOUAenco5v345edXiUTFhq+DBu20IrDaMeK5TURJ3SKzYy/M
JjuJqQrIgOL0lW9YmOgOONDLwY1ujMiEsL1rAOIQvgEYTNUt619Nvuin3ETh9FGcn0lf3E/aXLrR
QJg+kBgbjtnmy/Tpa+E/NsImF0KJsA/88E85jPXqPiPg44CT5v3ABQVRy9//5k1ZeKJzJOhCJAWb
EQckPuGGSoLVVqweQoqCPIYsrFz/Yrr8Kd/DtGkaMo08ifGaGfXrPDPGzs2h3qjT+ZWJQRiAD9Or
QtYr+kp0EujsjfoiPFnEpRgYvqF4yQatxcjY0lE1HOr76/HKiFIM3RUkIhbgnP/AnIlenztkg/mS
O7P3VYKiZ5FgfScXg733R8EReY8XOesGuqcZMEaupK9W5NhcnysqVFhlQIjm0hg0BGIBsJpVOZ4m
ZUR9Jh4jBPTWgj9GRtOWx13bpMUnMNgCxFKVx5fDbYNDMTHoC15/tk/2K52j5xuOyLHeih50Xrxw
X3oVuMYWWWHmO5btUh/4sIOJVQ76PXvSJfMS/f2ywelinMxDM4o8Rt0TI7Ooquva7WlFDcp0IRYn
igUegiKxNLaLkVC8a04pEs3SsacJ7J2h8KAfsn+TwSq7gZ0tZPMfrr1xZkOYgxoanX0pD2S6z8Jh
uugfftefTRrFZrJiU4PToZhhjThZxY7AwtFp9Mh4oahGDFS85Jv2tf0wjBRF3ycbXsOaYKyul/H2
rqZO9VMPkNio9DjJqAs4lXQeuvYpyh2kNBV4xPsRDdIMiwmmWAvqvP/ZXx+klszAEYn0l+KxHMar
s8RHqeBrHcFa8Al4hfl/0+sQ5JIz1WnkH8Zqm7gNDfvD5v0tmSaRW+9go0NUUvxYpeVIvbFf/1fA
yYKVIgmFyEBYmLpgAv20ZkkEMtmJhE3g+acPn9KNIx218D/T49NKw10supmHItUA700x+GSMSrmz
pX3FmxDfgbKmfxVBQxipqFLSQIuoqbAXSSlw50clOpXmpUwfQmYp605WBygsAsAByr+P1L4uCGok
4ZjtjqETQ1uk/CE0kBhZNnIyS12LeQBmXPb6eGX3rn9W56X6wffoLwQmM3AqDBuUklUs/OKgmaVr
v03MsX17ZCNmGJTSGH1pbXGDdv5wNstpOCZnYaYFAKF0KS1P55GabPRRe3R+L/7IzoaMX1PXncxE
IpBRv0XNN3EWE2goUQ8gnmNHgkhMdZ9LIZKcThTQ+Oe9dYUFarLKSfRdAwbhLdxzYBxxRPQnOc12
vtKaVlp9Dcm8lzdr8Q4ErDzHX4eazHEH4Xqqzzt1LGDKh3jCYbr+fJURzOtI+lBmFvQEow6ltRSF
0a+LMkPzW+yOyvYPaIVyZ18nCqixWWX6bn1SgB4GINdujc2xHKGRglcdU07dOPpgCXIms4eNH+Mz
F6shjNzlI8I33lNdYwD9eR+DylE5fr2txdDsnyUGyf3C5sej663qtcccguoALQ/pkGHnimzHVPpE
a7WmaUu1lBsjc7sPa1oBao173vQowSNapwbxQFy6ejviXLwye0HyknPX4YRYnA1d+IdFvxSqH5Wt
9Cvya9ronal12BMGCi2QoXQJ2ofjpuZZe/FYEnvlVAQbKWCLq88BgSxGjiKsY1dAmUVvY0mB6beE
nITF4zsWaOfzswcxUmmh0+DnmG4nifhmXd/8AYhH6biBrEwXPS5NblX9VwHyQCQCfn8cAcfILcgo
D1218rtTApI4ktQaa2Sl20RVtYjGJgolIILft3lkb/DlVTCPrpvP6tvSct8STZ5cAnwGldQzgDTu
HwUf2X+BtgvADO6qsYVIJ7aumWkt44crctjnUj7+RMpedKxbQ2mEAsYoKcGM5tt2O9FLEtOnYWwY
6MaUmFy9vTc2HKGevw2NNtbAIMlwAzJQT2qdXiKOVaYrqQuavmg0AgBlt+p90YtyuMjks0MnMnXd
hzFV9OQHYIy1CMD1D0BXovCKhr3inzyuTX0Vmw9XurIdFDV8TXqCQVi89JkfriHWVMU1QRNze/Q8
sOpIoAsS2wnGimQ8D/OfgIVq/KY6v6uB0c56pWVExdJ8fOL6dbThgxcZcf/hGIhWJjsSzdw1JTV6
zcwRAdF/S//1UCv2GtEnLVNE/SsK+/VBeb3Takhx2zhOAenBuMuBa3eykqfGKWS+V1Oy4z0COMb8
Zxis5ChcLZDUWXROWokj0J/gOWc/ROkWoN2HOAk3jJzmuOOykFQhBPyGhCmpOPkXlOK0eeX+YUu5
wuDimbtwmo5omaYFxKiTk3dSxvkyc2C35Kr6XdOP2z6NKpLWO4ppwdYHXOP26bFnuv7UWgMmXbBn
394f095uwotZaCFH+O2ZWOxktpb1mBy6q14kTX9jmm5iSFWk8bY5YYqCQ55oipkLk7mJwI3lyYHd
f9zaVd3JH9Wy0kND966GwSENvqJMB+yTy63ol+XcnEajK9YPMhCLA6fGSb1dlm8nAsQRpmpxWqXK
NFWcj/loS1ZBmwN+QDcWRFnWzhzHeTShU4ObHIgluyPgGVSHU+d1uKQaiw2qqN6//0Kw1gH/kRI2
cMD7VqeBE1mToVyS0KSpu1iK/LSMu/iHdRnjIW+Gk4jGdFRDIzQAMEhm7cAlfMCtdYRulrc3OO+u
hbuAKn4RqCqTgmMtauN13jidlbGRX+RXKQhRtzXNB2tDPAfKIJDgd19J9ok4rmX9QSEd3XcHlcsa
BPhnepnT9aPNsPeUkQKOuUCMJmPVg2HlLtFqwq1wJP1j42LrNWDHjzo/5k8NrbaOjitKuk6m0elK
If5WtqOCOQO4PBYYPqYJpyzuNS61vgSTCwgzoaW8PJzhHSe+Jz3XzTX5Wjw1afYIhb+n44O3eytg
Nw0t/RF+SRtLrtAf6KZZ/X1KXqJhC2LUSDU55Hh5wA7pt3DzyYNgTgL9WS5FCmPNMu9tTci5pXuI
BARWLArevoZR1y/BNGpIJsl+IlfMqegKvKJWsGrsC3QK+CbErXkh56QdlF7Kia1X5GOGS5ywasPo
FmkfHSKPIEEffenPAK8D64w6k66KVs1dN4GBtMcb4BV94SB3b4PfUFxNCX83HYHDsXR/MchyZQCr
mvPcaBrwDMtZNCEnp4z2Tr2QNvo4Nh3C0ytKL6dJwE40Q9WPKaZM8tCANNeBXLhsDCFsFNnznRCK
FJA4KkPQFTZaTvOUf3plHw5Lz3RrWy3Kp8HXsWeU+erwVNoOpk4QcZxmE/XgL7yRGwVWkPg9R4kc
UkIsOrksmijdr5ZWuHD4otd2cZDRJs10x3Mdcs6Sqsk3gKD4qJ7p3as3D8EIUJUdjKWUS1AmsOAw
tX+YVcoSd8nmhXC1444PGtX2mkR0RkGEULVDGGG8IFxrHMNQk6u3emjJlek9648ADg0UWdjtLLEX
PJqJ2pqpjNu3Dep0TrAVh/HpiD3YretwxtEsqHk1JOhrGp93SivMtmVSBQgM6iiV6uj6gX5Qg5AY
49jrpXVJqSfwk0UL5+HXf71+0AhKWG5+qlsrT+/brlO0lG0C+kp2tRoUueiyRp8jjyK4CWU9gWfQ
soHkCh6TbJfsEMQErVs4v8HtYM1DAbARJ+qHHTkv3Td5GEJvkwEznupMc9fh94WbB0BLqdI70M82
XilCe4N9luGTlHHl5zvVSc7bFYH+5i3f6XbM8QeptvWGWmztBE7ujYowTMCIT3XVBR2IRwvewUbW
LesirvfG+rWsg9KCuTxu6W69tzCCzUWqR4QmPT2v5S++i1OmsjIQng4pWuShL734Wem+gTfPndJF
Jbxen6uYgNzF2PNpBgNJuWGJnar3WtkCoUNfri1KJAsvKPiZ4jyW+Eg4tyA0H27YGPq71zd6iDeb
/sl7SwCtLBvavqKu1RMXSntHpMzhP89xbS989qTag3IGShW8pY9lfR9cetnjuXdkHQjouU6a4Etj
tPLfCtITKdHVrXrQjVD1hqjbSiuYUX8DJ/g1R9WEng29xQIZ2n2oTuP46s6Vml7D+Nja2OdmMdTP
HeYTY20Ym0rNaKV1zSwRJiJuKxxQnBu1pd7eQEHcUQNOKWAf27C34H+3TVYJ8NBPJkpZu1LH1ql5
bTxOqgQSAEy4XN+iI2eVpTzh4lOp/Rfddtt7IbZSVKv/DJPKTngwu4FHj75xr0GfxTl7Er9aEftC
LVBQPAzdtin0NIy3WmwGud77Xyy3THto8AwrF4I5wjiCUYZliaa5FpgTzsZRVevG3AJfzznzMqDf
q7Tfac5M46Bo7PrgK03xV1hO9Oqo+HcOMI2j9Uo9f83dXx4TBdIUsI8H76s5IXNV7iZ0hIbAYZ+V
YL/pOZmY6xK3T9mXrY6HgKy8/T9xaH7f6FFM6Qo30rea06gFhZYngFOaX1iyJPmWFq2Pqai5ra3F
bRqR/y5cUtLZAbsizdJEbPEYOyhrpPJzmcrKSambjFrP4v6gFxK1ctc6op1GQcUNrx9Ud1XxzzN2
zCZXZ6NrpN7Jt1MLqu+eal9EnBxBahkY2VtNe9sRpizbUHorUhMaD6cvtOhMqo0c7eOONfB+qti2
Eu/0QWeBTb9WTbKvcWWFfO/jP8pizLiYn/kThV1pSPutIJijte+eZeETT2SFSaNt56tweAOhW7l1
foubV9FeAZW/1WIBGJdBT8QAH9Jjonepi4LNEGPC627rapib0UDSL+LhfyGCnM6b3xnGDfujRGmf
KlisYz2zm89izIT58FwVqvYTjgrTGRKU0IjBuqIA9dIzW2sL5s3fLbhFBrZRF0C/vSTuH2jpHz0K
XatDEbZh3Gd5sD702GC8t5uGbvjwsxchdk21oG6ayzl3MW+Oa/hrbWxgqA7EFp8UX4/1erQmbj59
Pu2d37BskwdpJ3jJNGZzDwiLuU+kn/QJ0gmbuZVH2PzEpYQAuMuuFN5/3D8TWhtiNYo3SIPzuEwG
h6RogWu9Uo1gJow+L4Wy10KmDdRFPICHV6DgNLDZL4S68bhRdmXNeuvXkv+YrexUOI4kDAQIpwnx
8AqPeEeRGaQvgu9cCTueNK3nHbPgcOSvlOOxkdLXte54KT2kARzsokSDMTSDibrwJlQnzdNW/aaE
JJkNGSYxpsiUrkNjK0/EWXVSqsrmux78QqaFr6wCJjVPK+dvDaDBgSruAVEs7vO1yIQDAR/IlLlQ
f6iLh6HdKXqw2/k4Z7/d+ubHccZ4vN4OCGaGKAQl9v+dJNn1DvlsQxnVvJNMzc2bPARE+IC8KtcK
U2e7Juq6c9HvIaQ/CLaMI/7LXhylYk+BAR6/iJjY39etC/PR4Z1d1dDevuIc4zx+2cZN0LCC/07v
03rLmfjUNUs1YjsbpRMzVTjjiQ1TGrpBHpT2Lp8GfloGQODW+xhj9h526bP0+vj+CLOJM4iSj+qx
MAxDyNM9X1kYCHado/AvFsSUsMI7iusvJUwxf80MBGGSzYHK+pK1zjgS4o084Z2BWC5y9fxV+TZ0
37c5HaETcU8kpvef1Omw8SNe5JTlcrfdtsxkO1QqDBCt5PGwkKGysi6uizBFHgTHNotMjjPNOGB7
KweU2NwwddrsdxLDgpUqjffvzgAP9tih5a3YsivQ27RQpu0hQ6iVCpR6TdTFcNpL7ahtX4ELW2O9
xSWMWL+AIecYo19cI2R2DjATaAzXBR+yz+vVyiTkTcCsIlSWWSvRWcc6LT18orWZSNA8vreN4eN6
LR2E8vMQZ6fhGM0ClPDAipL0OUn+zszT7t5UpUgEqFi5pGnDsauvUc+DLKZ0laGzW2+NUK6UzgE2
gK34HGoAuOvaDYq3EFVUEWU6FCh3iPYlr1JmPzRNB6pBymqHhD0T0Yv0Zi0smISrd3fYS6YpGQO8
cINTf4OquY7QpU0wsU2IrBjRBOCOs78Bvsvd/RGZ9gNYP2sgV2Z36DVjFfq/C6E8vclMHxg3D/In
Ty/4nseS2mMOq7PypadL9lt5/wfh+l7c5AX0Z1Qfdt1ZFxOFCmN1jo3wx27gOCeaxn657QyaRJ3V
HQzPqYIRKEHGOE+xqOn3R+brL7lSCGP4OOJ4ndVd+ly5Ojv8mndvjczjDDbITFTKZR4YD8e/E3Ws
LGsS1ihm/4ouAf9V/VgI5H7yuX0YJfQPex5ok6X+1HTKW6vNbT2jYwWlOnmUXywhr1uMOHBltvmy
MBPyTupiB6gDVVGYjl+onU6jZ+Lkg1mTTnR9bSR8+XZd2Z+kQNs3TWiiRTSIDz4PjVOv75GSRm26
tRQU2aaGkC5NB/PaIkijJG/7AQeD7Vu+48ptmOPI3AeD4cvwv2jPSscEVDwoMDPan8SDxfSAXMgz
diztIxP6KXVg2WXdk1wGmkiQLGgNk0R0PeBuu8j8q4gX9CvYRkAIE9Gc1H81tVl32Y7Wx/ZUkx7c
ihm1oro2JVrgEjyMDJk33m8+PL7Ib1u71d46gJo3sMoydqnib11Z19S4wk2Il6xgEAfgo2SRjxNR
h3NmsnL2VY1ugsGCy8mFd3emWx1R/Do0rXwz/hJTH45nSldGqO9EL7iXHCajThwICbhWKHgHnTeo
t/1ECUB2yzYFbT2ikynA83Rmw+rRuNCcih6Zu1wye1A1iGwbdotlTMH9xg/3mzFsAzXu631c0t10
ZXATg6wLh6fyCsbh5Y6k5oDZqhvBtIfuWJ80de42wyM6M8eZJu5jCrvLZMA3K5R7tXdWgTywcKvH
d+MrFm9b3N8dUJLkw56Glf6hlq5MqKTfU4O2RU2LKhs7/waLoWM8dQOOv09Ud/vh1VMM6sclGrGW
aXqbg+nA2Mb2pdh5If8m6lZPRHvc7ttMlIm3LEi74GAxYOOnRVG7lU8rR+Hb94xcbC5FEN6m9b0S
PhjydNeHuhutfCJi2LvMfCsQPjbZKbj4k2lfFU+pzz8zMIK68LB2vY1ci3tQODaCmvDxZ+TTlVSh
tOSe4SGoAkYCOp6xEXmK+8ap5JR7Q6rMTf8kQu55HRBP5HSIM/a+5Z0XsQaA5Qv6EWr1EJL8ZF5c
CAR/yoUnsAX1l3hV3jMdmJiReS4gJvNWqaU/FW5YJYe4CfdONiDQ84dNpa4C0aK4JWCmcaArSJZT
wRjpTf6fRvGMCBpzGF+EQuIVLandpKnyBEVN+Yd4UigOHc1Kl4i2cq+udN65Y7LOsFfCZHjmto0o
jXVtbwNPn0lzGpBSpR3dUyestwb9338JlnG/7cjjFVI8lYCsyJPQqkc2CGIVkRlDNxhuV+7ikVJz
mfBX8lmm/qQpGUn9PXE4iFkSXAgwpkh8hHYRjqhskrfgZL5RsHgi3KoBY1+R4T+7p817LvK7reUk
IXsMLOlrKg95k0allt23Z4zdwzjTdykXDwaROOgfZ/qqBEYtyEqyorLmwI8HklvOcCHETmp/LN6S
JFh/g4y18c5Q7BxVh4ju14KwqvGHSv81HXJBIKqO9iINllJ22PSposzOO8SXPg6FDf1LVHZkuY4z
zNMkWiB3gdNuSflJUJPyTupDrX3BYot93am8aGrlQtPdmgqqNJz9eF/5V9mFTi+45R/aV/v1LTOr
/pbHPWqXnT/PGuCg8xaOLFDPxe29hKVr3/D0I2lUyql3hfldJqZstXrKxOG6woRz13PsOPSeJP42
RDETUWj5qvSXHWNSWoDFz09IirnRG0S+5fKgSb8n9fJX40CLqNTQ7P0g2GRIk4kJFiEJHReh3nm7
rYQLp/bsdjbnD+0PwjRIqg4UuqSY6c6jaBExh4LkYVC+57iHwYKm4jlnWIUVcSPjXx7sTnJT7SPg
Ad3N+WCCioVHHMbFns2FYi+3Zb4gEFtiQRp5rVxTUQYLrEXQrvPj2L/vwXGhmAyYWRs88ArNHXNT
Sram+pPcWmhmgfN3ZWSkkw+EUo98kjLbLx0ZlQ6WWam31kjHCRNl2pq2OM4RVqrtVihDo+h5i9GD
ZmnfxxkDLmfdHuFWmoukFQF4Z00fNHOMSGCZXUT5CQN/YT9+FkPCQNHlTouulMJVpU2ONAQwAfn+
nhnQI2mWw+rEpIRgn2C64Lk1sGg6f1iWUdLitWJm4tANIWpsNHVJ1+QK34KCQZEFSm2bt0k74Ot9
81YLlQ7ZjkkKmudC0YgTm028UWM13u+MqaiMis0wyGuOfjhjdTUecb2BJJ68n12n44mjeYmYCqFY
hBsDQ6oC+CqA3Oatp5YoKafkPqG4dUQIlzYqEvgdP49GsRYofkBrSL7LwoHyc8eKJJzVEYmuMtOm
UqqRgAmgycL8Ag0oOWennVXdfipOxHiqSgPyjE21nkzDM5hD4jXALdZMIBYswYLEqCsKm2GKjHmJ
zRA1NHC3GlPHrFBexkP9CMiv4ZxKK5sMiqbbBHIGh+nUlud3ARvcUo3wTIyaMLrButdmRYeLHYE4
mWkv73ic/Ovev7uhSu46B2gSAH0AUMQFHmbyfrS4WHYvGcF7dXyxCea9YDOBuXHJtQbYE8IAQtMq
FNeFH5GEcY7DS+vrmHwAq7Nvdc3QgjDt+8w/RML5CNM9XwTnBRCpSXdpy5UuX+f4d+/QcgezCpiE
bEeC6MpUaMMfEJaTRinGXO+omZPeFqxOFwycdWFRQiC2aEGell1atX6HuP07215+Bf3ft/t+6cpV
gJJe+DwlaoN9K/cmYdtbudfuLTJpRgXw+PqCgCWxl+eDrhvyKO64e8gsuBjeTQPQF8md7BaesOkR
MrUXFIMuaSyMdjYXRUcP6kYeOrpOtzYNcCKqW/JaK+2aBXrafL5vobgybrxUbRvYMZynEzRJFoVk
n8eEym9PThBDUADm7sKgQj7AYwDGbWoImaHVliaMrKWuURFfd1TrmKpLqCREncmscZUDls32s1mu
DfRwT/2INOo1+v66kKdK3ODITsfDMD7s1Go4gRtwsi4vhB6EWEiNs9ECiJfbRoywPFeiY8OwrOmh
uMsH4bteAqb0rZmrv8nuimkXXMu/+9h95NFA8y9y3es55q0gkU5YbepES24dbVa0rwiEM1nlxBzD
kv1C7Hx1PaZ2TzI8WZERf+j5i4SZQNAaHapzfFwWIG087/A/Ae1dJkl7feZk9zliGG580itgmQx0
csLZNOJICG7+S+sKi2nq35F2URov+rXECFYDDok3y3Fvn3zrhdwLujXY0ASeraYi32dAepBQtos4
ypyzE+/S8Vjm2CGC4WARKjjMilbjyDGw2hTaOCNfbQ8iyfSKE3a9K5xRilckp06tTEErQn/oTX+j
WqMpCzYYNKGfX8rJEziDXBa7042IhL1lOngLjwPEQTmN9RcCAuloRtyrCwXE/I+Cg5N+CAT8h7iF
zU88dFJc6dl1zv44Ulby+/2injLRRYfkIcLYS/eKA5zPrJqABVV59ZL6SoBWpGQJ/FP+6jOGhC4I
9y4IPKlULA2ypwpq74MVJZH3UzWKIbTIIjQ2BB7MGkqAVEHCJ916fADEHxLqt2ZcRG2zdZ0hpZv/
47zVPQbgAXgsH8Jbhpa8+Jn9FUpiiimHHswEIhXOGXdR55j1eD31mQwgOso/cSd0sx9kMn17HEDB
kFJQTuKLBHd9J80y1Cr3h02Vg+q/l9nXVPr3so4BAgEZA8MFLTfjCUAdLAOZXEtCZhtmjhxwZVcn
611eMajDw8ogCZywjc8KnR1XK6KZl2tRhyEow52i3CiZ4Rv64rUmK+vRNKrhOIe4nc7FEytr7+zo
hk4yEuiU9YYdLQ1IYfupXSQD7trbvPcI4/PrxOu/+rA4IfBR83Oh0NrsW4eayZ5MdQvHwIIGqjZL
aUu61ejSwaVTqJYDiTDfXdi2h18ZylLo+OVaqAC7U0aECRdqflSf2k1nkxh3VL4hTXvlPw75ywcc
QeTd125Cc7Y9Du5ITrettDGg4bVCVv3p4qae6m4ZQEW7ukYzOVRojmRfCejmEFZStgHIMS/TjUni
M6gQDroyjfqUmBSzdgd9xTe4w07PP2VNcgJipC59bTB1LAi7wbJkmC3X84ZWaAFzTzrjCcfxNli+
Pgg83VTNQFpqwnZBONz5E66TllihUSfaCKSr5lyjnIarMY2EIFT1q/6mKo0jdVcenjEgoOa/Z3sE
H64S8JBD29++MOA+gFUWZ8LHjnJRJClof22JIJ6IZ1W28A2TfsxhQ81Wi30HK/Xh9Z8S2aPmtIr/
CQRSStlNjX1QZGhO2oVTIwfNESqa1X2YCU5yXwFSByTT2pDyHW/9eq4vWDHYw6c2+ysQPtMkr6bL
AroDd2LDKVz96IzHh8Gj7txldGdLvLelyvk8irIZRyO+aKgdKCpz1MI4yrR3O83ExfJvBvsX2W+T
2YRs0ibhcZNMC9JoQ1omqkjUfgHsL60G3ec2X6rpOTzxO2Ba2SwQ0i/06T+C8KhaOmojz+qR6Ldq
Mcxb6oLtFr/aanC1GoMYRZhr3K5NKIF+2maCl/UmigBV5on4uklGWINEJYCcNAG6hWQ9OIKrBqz+
eOwhmPE/Kvpc0b3RJZqluYVhhPW6Cov36HaVAX318+t0i8r9PpAFOX6RWFlZpnfVG4r5ey5X3Pmj
S8CdouKSOSUAWE9u6cRqoZxKNu4WY9khHIALsVB1ECP8EJ7G0oc5b4CaXnx4d/zG2aS45VGTFyT0
vWxfmVApSZwra4IBdiJXt+V8cjyUzQeMMotv2jmJT61YEF3dqcESHdwCgVvmTSxJzS4BkTgFW5x2
qkJbsEzshOmXHxA6xmoh46puvvq+dmLkvpjOPbRV18szFN7STh2D12MzOyR5Ua5POWzRp9x4+Z9O
IVuTIym7seKsvBZA3mZ2i/EJcEa3pVYZoFd6VK5sPp3eLetnHEkhlDKo1ZTG4/OCCqUSzixvnORj
4S1rbVXDYSYFZ9rpGW9WUGLfkKM+qkVAL27Vp3jXskmMF60SPFezOHc5Rj4ySB3DlcRWljLcdP5a
Yd1dKsUN0magPVsZwZkYQVDFfcezras+ro08EVFLJfPNW0V0x1filkjDWz61niEz7y6B9e1RCcGJ
Fr0sCTT5DEQY+0JbVD1BOKFKbrTxcN0a0PxFMBikVQy+/crLrQ+46ikrI40bqXBYjhUWbSqSCBHx
jdzKA2PxYvfJFKrlKzugQAUpqNFa7K9N9MwGyKYqMt37pVMEvJVaSoy0pcOuWYalHC+7yFRB/IFE
cajDAfCtigp31jZTK9EoPFKam1pfiJSkRZpuU1rkjpG6vw2luySPj6UoDGhZzBRGDLa0unmYmOXc
OcTQmAbASlKFK9xyOIdXEKDwTiADyx0PJpafmcaxWMH0q8wse8fg6KdT4BefklI+oDuOrpyAV1H+
agCLmAQWjJudkh8vpghlJubPVn9JnwcAHv4Oo6GBeV9BHbpdbbhIMS4GvxTBDc59f6xyC65Uj3yc
SebtmuRwCc3AG9Yn1qFUcuCBKgV2m+GjwAumAJ0ujc4KVqalDmryHagKOJlMqpVfBQnyj2QIpGrW
ACE8EDFoDo6Td1yqbKJfKPp610HhRQezpgSOMChNnBBYGsjjR0RW2maBv7awlkWZ4Q8UwEyjOjs0
DoThzGQXJD7Mtjzoe4CC6cdMUvI1LTTjUp6N3+wMS5Suj3NEy5M+4SS63DaUE9jLM9oVGFzzXFFJ
xKZKK8H5KtclL2hKdGAkaGBmJNXmdqlvjf9g9LbvuoNXzMNWedBysRWZjK5iVYWg/BhpxAC5ccZq
VBWmqhqL7CcfqCH1qAXbuDBDYbJWsYgSSZU6nFxuU9qP3s3lHyg9w351oOB9dIj1ZAQFU0CizrVK
LvprwhtJtY8NzjqADpF+iv7DRqzxY1zoIqTbaiQtbEWgrWxXN/zzKtEEdLQJcHfOd+8UCay+QWuh
QD6Fxhbaj4yqm+X6ve84NGMTQSx71U8hObfN/6Id6/5cSrZ/9XiY+wcRpiMyAct3H1Lm4vt94tbC
psnv5VJkM12/fDlzCIYqOGz4EbpOU59xdVxBO32y5GThijtbtd++SCtvncSjFChrUgvRS91idsjO
YImft3Ef3SSL2NJUHTWVnWMPcBeAlFFfFWPiyb0H/Rp+GWC5E0qHQCuJ4Sd6awvxpIIqG+oh40Lk
e6N+3vJZ7tsCnIBnglJ4qT/3Ei5KF1tj0RJ2szMogpwvbqXLHHs3K/XA3zx4VMq8EMa2eitX+0sN
8d8Pfl6cD2FgDluie7RakWxRxVdbF5p8KCohdd25W1zSLrFS6IYW267DwxqhWKEikIjvlNqLzkZE
tZ42D5+dS1+CFNOgU3M0BTemvV8Nt+s2wdbAxQ5aA24qqmVpGxwxUUxr4jKMblMLQWf1k4HWStCq
Wi9a0D5iB1+YNXjbW1nWjkhlxDfnip9LNA/iq4sgH1xL5cPWLWksf62+6KdYyNdajxiFQMBXw7M7
gxkwSaacms1JMbIv4xJ8HF8gP6QbEdaQUmyr1KVM9aNbvxAisqKQYKtZOtK7CL0hPEEhZxFLBW8i
Fdaj4etMZ+OjniYYIjNy1T4kdJaq6/ivR4vSWi3U7NMyzzQrFwWceTqIJg9WJJsNZNX52T2XD02A
tc/GyHaABuUy+ViOzV+oktyeYODLkpNjrpRkwUMY+VGIlfFDfm7UTdRhCHA29k5FOEfJWyvGOHuA
73VyPSZgmbD5OMIksnWl4AcS0Qapo8bbSra4jc6azp/rD7jxODw58/KaPaHKG94yJcp7Rx6O123Y
YHLKzXVwg4vCenSXpX4R+gcqMKbfKbxVKfOhfh9bXO4pvq7SB1fHLQ9IQiN1MIvBVS71utS78Q0p
Y7WhChP8P9lidU9QcvYl66HdAT+qLTfzaq4n76SVeUYQ6Nobc6eZ+D6gNMOqqpi95s0iCZQ2Ie+l
/diasOW1yWtCY3BAWhh6A/0U/cB2g2KUBIqGhYq1A982bNTBwbC6sn7+lc9xEf3GAzFri1DR66te
UcapwQMfZs/C9ByksMJ4UTd9SS/zECRrFYRl9IHqXt3giBTprI846cGa9KzRr8uGCEnhvWd+uGYi
Ra2DXYRHWJSKxu6xX7pmi4JAGvkQ79VtxvxD8A9Fs/4lScWGmauy1RP8pArLjgIOmxG8LzyNXNlw
mO8xovq6abzqo8xwwuJbeDJ+UNyiqswK+VWgJ1xzyjve9/tpuhXRBBGGf9PM8IiCQBGK3RBlvZE1
j3eZ4zeTAB5B9cepqOdibmtwtA/pECQp112ahtD6xgEDd99rDG6vVK9Co8O2zCVsckiIThS8Dzjj
/3tpujSLPfzpBiHwEjLu51Pgap68mgGq39NO3eLC2iUTqbVsK6VB5dfgQKmbjJpqU0qX3YdAGvkA
8KTW3fj/LvlRkjdhcYnJME5H918yJ6O/DuQfLS4sQW5vLfLlvsSXfcwENsI/6pr7lVvyKJHBWmLc
OjjDlhATOEhztIAkd+lcLTDyJ9w/PjSIKqX60VfyKLIVt74v6zAo6IP6jZAogqtunuXNXVcw9KV9
RokRxkeS3uzKtAVntLmTVwkckoFemO5WW1nsswSrwgCdA3/l4NzQ1exgW3yClwbf122+TEr93tBi
CAOmeerMA8z/b48TJw5dCYpnjI/w9YwvkQO2U0WueAW8H41wuhOJVrVGFKnmLCYwKJpjUQWmu64m
vvSeyEWojRTCTtrszzZ3zAWQhR+QwueKCFElWr4LfI5h+z/SdiCjNB9AS/JtFEpHvMLzA8oc23+Q
SFJDz7h9QURe0MxnyYbw0ZkxJ7+fAXV47+9/65znci/ViMDkzpOZoHPVhnpOPzAr7ZOuFYje+DU8
aeyWwUEg4qML3SjYDZxIqdWNKsf4AnTIk05WqKiMKTaTgr4dhPdvCzBFMQen47s/D8gSXsTQnsTG
c4cwQUwgfix6PH3Lg+8PoDzFLQTJpEVRcc1tbkIt1VXP+HX0Cz5u4IFVArUmHGu9xowyD80uzt48
tVLrp6GxqnCn1XmX9PAoJmWfDYEbayUKPPobTDRUuC9tsMECjVtgcLgdD6pFOltKNhZQBC8l33Ic
VrMt1S3FzpT3L0bBcavDMP/e/hUs+8gmXTouG9yBthiOyXvDq8DLsrWo57GlnWsaBLhBX/wv6ipP
sNELELtGIpFpHcUtdMc8zl6PCbDQfeMO3FLibvdZwgbclgpFSMwTsuHvZ2bEonrfsqb7jGZPP+gr
7CDw7Qy4yxaZNwGMgJmnGDHWRuhy/Qshc4GONcAMtO3o1OeNRVEAdCljJw5tp5rx9TFcG+Wu7z1H
6JA9xWvORz2ANbcMeQyhd6VXRwjtX4jFjlL5sfHCT3A16oyI4Z3geC/Z36BUb21LNITxNJYxBVe4
QZ2tT6ODQfPnHG28m2dyW47qh46QxaXX43ueg9kfXbVcv4DG+3S4Rj5ceFiVCOu2RTKGW7Leoc4k
V3YhOGFn2RDWtTx2ftPwVkNdBmyAWpvCaUmnFtCy+B04JkuAMl/9xiullm/EzibNdt5x5brlj8Rs
YMySLlyryijiR2UajHuqLBh2gJUSQuF/Af+ILVdwPKmXTSkjqiljYNDrVlmShVLJihL5HSX832ln
fBYsBZsB5ng5qg7TAYZlFmYzvAbfykUIEdkCHieFuxWGYvTWOUpIOQTlgbno6U4kpm2NX4ReEcF8
p1UjTzrLLUEcVvVtc1UssrnE2HxsZp6tvN7xDHonMnJR7CYk9PRDahxBaI7zlkIjRpHph/Ei4NN/
NmnjOZrhEtsQgsUx4/5MvBQ6gfHn0D4NypDS9uYZraxdpMTGtzP+RUxoXeuHJ/0UkQgGx7RO3diL
R1lX9GalENqfFrtn4W+joH5h6dtOPyNt8FZzjDPIOw9HWdNPtKFYwrS2vFN/77pmFuYIxHXJNtkU
aTXDfFRJKzgVspsi6qA09mSCu/DkcWZagOUjFTB/RTkDULtW3zoG7oPgheLdrOqugY5eGK8P5ozu
Fwn7hvwpAHXzHGDm08AyxS9+Q9CQ6ahsNqjH6ILo43+sTRvh45Wsz8GdEzFqHximSp652EEGU3fv
JnOrgC/q3ddzHoZX5ZAUa1JBXKXjwt2z7AGrfGHHbexsi57Slnky1rXZrC5jdTFV/dIfNcUbMgYn
qD6F12EmnqYkcYeP7fl63V7QQ6jUkJglGDGtC0GDsjZwFqOAELhACAwLRveuw5CA5raBT6BgCU+G
1cBH/z2kbDp45LJ7U3U1PCOOBR8mbhxN+XuQNjxsuPoYh4eCRS9V4f1LURlnjnZazaoiq/w0OG4U
qvdbgFfGPbnEPqoZSirKC+Drg3g1Hzr3TDJbq3OqGWkg3KeMjYI55CJSdR0B8e4maSi7bgLRkr5l
yPsPZ2IPiZ+GvrUpUequ2v6SoJvOjlroU6Tq1FqDkMCCPKCSKdHOFsyJqouqVIRPdK38/R6jhIIH
+UYhqstxT0OLkBLtNYSLOW+MAreA3qnsZQt+QDzwyYmw8sB8dV4HFOnlZoRWqNYtQ3FvJE30aTy0
JBiWpFJ8wfItsnIfg6nkK51sSuQ+sCEHP2bNGHVe0oNcZTri7vyjYVJ7n3xM7WIrwWReaYM9MY8W
sEtWudzTjcmvb5WK3h8ucYgnSel+EJH8qLbTz2d/TzERoo4ZVeNqbTL1th2Q4RZS9tnxvmryT14U
sgaWeOMLeVy1m8D29OKzcvqAdzQogJIIt4BvEiu5zRyJD7lG9SgRQI6wLgr1EJA96IXxFpTqWMgQ
MmerHoYzARO/ODTakPYj221zmeKrANe1WyjDR12jvSh6lNYWfpGKks5LtOAtQAWGTkXv7zBaR34Y
DSQ0IFvGlTDvn1iuVB8CYHbPyInWSYw/uSR6VOKVjPp0GYeCKN/iwtOkl5i81RUiqWpKyJ0juY91
OIAVRg45g2qwTvVmtHOANe8ymjhEzKuqr+N/3EpuuIAi6bciBa61NY9Ad47vVsndspxvVpZnITHn
LY/MdPjsvTdD4NtvJovDki4P59ys4nwLx+tohRL+QtLsD0b3Spd5+o1AuOIyynj9oEZ5ItGpojaT
bfT8JU/hI4tsmUl/XMVi75QfvGbyIZhAiW3jUnObAc1Oci4RH6YCv/5DY0lcZsyzpROqXs77Zn1n
lgvBuOwJAK+DcP/xfjUwyfGbptTCOVwcMG1/w/1uqkKwnJqYVDlA3jZuE2+MZ67ifgntmuP7N9x2
gplto/SNxiFTjB0ZghI8+dQGg+SbtDICXyYlfa3q5UtrXrGYz0DeMumfRECqa8ZE5dGCusy9t6pQ
7kC4wAeCAMsaYzn5XJYbOxOdeDLBDRLiR9BI4eG3M5Juej7fIrm4Fn9VgLJYnLEXIK53M8OgcfgF
Rz/6IQ/fUVkr7chmtOGWOtrkX29zFH438/H3i+F0+LWMJEgB+38Mz1vv3+d3xJ+wb5htvWu25nBd
IOXXfkEnQysDkW41f8heQkNx9tZvg5NNPi1I3BwA0jHwjUgdGtJ52dl2ZPK1PBDFcO7DYkhPTe1D
oJMkEll9IeSCBlIabE38M3UrF55mIaoaiOwuPKFUD18UQbpu7JqXh2khi9/j28LaGvmd3v4DMUxW
682TmjGWtBI3aKdHaqISL5rLzrn7IV5PrSIlhr+ud9uKkxiFnMgNnMiHX15aqmwXgpgQyLxN/V1d
WGd9c/APpF3g0hV0JbCxKnE5gZQEfy2nc4XR4er+uC21H2iaYzjKZlJBXtx8kDJUQmpaT1HOrC3i
/qzcAVOZ/ij3dIU7cnW2RsLHLDnSJZJrsJdhujI5lmGLVWdNuUPmYTM1+FtMEQyEibgEzEVXZ+37
7E+6t2+jce8BBi4A3hctU2N9tswee5qmaZ6bzBwgv4c3y/YXvxLU1O35BXRfsyMfUMnuSm5dKfGt
gUqK8IJTeHsVwMpCtxM6uYaRXvkCfzuadeBWojawBUWx3RH0LG3aYr73ATGxwSXYf/6E+SvCwxRv
ICaGMZuqsPZg82Qb82+qlFyKgYkNJ6iqkWdMZkDqWHHeJ3q+FsMGjJ+D2Ec6Z0IlKcKa2TqV/ec6
y01tQR3cOL0rP8Mzx0dhdc+1+tiEV7wDxdN+TDZUqrYlMffK5pdf2ry7CRDvmp+gvNUFNTWFlFJn
QsQ2ROQeYVJbysAcx2A5QEEVVucQz+qv6jTc57/COfl+OVPxvNgHfiTfEiQzhy0csQRuHQMpkw9x
GoxcM6etP6LmyRX15w4f+g1Nakpbm11tZIaF8Zf4MYjTnVg57MhSxMPFMWvzpUM8ESSlsz/L17gU
7btdNKs83ndnlTLVCjdXQmoe6ERipYvMSwor/XmXNHgCKR2/qmh5HpLcJjdzIe+GspzAJXLLUrCq
L4XNCkUSDH/FtwtDrKJenhosUeJWsrs8boYeDYK15BCBMPK3rcxrGlw3ZTtQrVS5hkoCXbFirY0U
yqHubm6JawKB4nZEdtNE1WDJkULlhyuOmFbtu9W6s+2jhI+aW//fONVLOvGQ3lTghloyrfHLk9HZ
5cx1QGt2CQtpDxoyS8l2QPnsLI/b5rew2MCUQmN/qPrDQzkFRwKEm5S+O7BwzOOa8azJkQKUWDkh
6MjKcuUdhxwjRYh/l/V8XAeA0jFblT61MhOws8pd3hnCyT0wl33XsJsfC7dMBjwSmfWKFAKEqQCI
o3X/Z16/Ofecd7PDXj2MxXq25XIWzzrXAiZsYCapdD+IhPp4Wg6QPHYo3/ax1DEvzPfIk/9RHBUV
GA7horSB3KAVqq81XsNl9oLVqsj9qdSlZjg8Ejz3E4uHePfJQak635j82IF6q/cl+Y85OeMU0WHs
0JaPXVG7Y9yaMpaE7J6eqyPJCZ9ySNRb/B/7pJJlGgfF5IUzd/DuUqP9/bHN9NPxwCp+2PVvmyP3
0oMDHQYrzDCWbwnb+54MuMYUDX6v7V1q1ZA3QVAv6MZnOrFvLYAoYFxEuN97YNjJSi6rOxKq45Gw
8/bwoveARpEFHOmRQpRIv0FgzjAEp5maJ020QtX2SJvSGza/vjjxWe19rRr8WvbnAozQyslurW2c
ZwRgagNuarOc5T1QYTkwNCkLA5X0qE09uqTSKcXM5zdqJEHsbox4lNiVYxcy8KTnOvhecLwjoz0B
df92xuYQEj4iql5JRZ0f1TkvkH/5vGWB+YwLHknno938CjraxweDuewyWwu8xFvBhRyYiY9ziQkI
xTpDV8iHUAsyL25nngyRlB/f9jEzvqspQnFNpZikPsB9GdtYQtcc49kjn4nmw9qGzDxFpfaGrHCQ
UMbPM39GAUrpb2PuMHq3zVvcmZC61q1s5wI9rDyQeaJK00XQ+DQEW2sVV65tU5qbCbMvx0zAoA6B
tCktWYzWo4rCcdj2D2JSxErOV4ll+Boa6gwgg99zC2JWUZTga3nBxlehK3FzHrP7YFMSu73GfBFz
kzSg6RrAdkqyvcNGx5WFDHcWUhDFoU2TYnVrEKydKidoXyrJbl3M540UnbGQECEch6EHKwQlL4nI
rH110gbg7IBrmULfMllT+9Wx728rDgpSmM9JNRw9ksnfQdMoWj3wqvTcpl0dTVvywG0pamOA/994
rKOahymcMdHsBw7gfTA43OqknjHUEIz7csmAR4o9jMA9UWhQxZfszfVtPlEu4pTGNqhz7qymdvv6
FEPIOiJ7LhYeaz/maRWuCLnYAsl1XhHUvmFvkYR6qsnp76/NyhjfLOrm3viUGMSaz8/j7Fo6KP+i
4IChDoV3JI5wQ0Cf7P6vKaZRDxtjj1v9p2VUO2g7BNo5R0YWynw72YaCR5kq+QU0kmb7aqAwY1gr
5PLJR24AMOCrtSKY1uEmF3vay+VKKghpPZVfgf4qFSuwlDBBjn6Iyf2kS0PRatZw2ya7hJusQ373
qkCA0Ovgpoa7Tz/OVnxxqLTJOk1+YuBLH0OcKyiBV2U7boL+HpjJ30MEF3S6QdXk9OWQLRE14CeZ
Gg9H/XbCiSbt0ToAj2NrZ5yPSUmysrslfRoeE2Zj3B6uS4A/m4bV/pNGi8GroFZrOgyMLtBC6atd
wl8ZQ0tGWHiF0dMVSKSDY8CRkOI5S2vBUGid58dVtLqKmnL6fXuDI3CskFH481oILiDqpC55joXl
IxOASAwJav4uCocb2mWrI9c/7ycq82pR9Cpt29HXp6zE9bSxMFLsA4VAGVv4EUPV5ifk3i1ALrPl
4TY3LxboBnpNBfXRdnGhvDC/2vZ9o7JSQKm0BvcasOdWsus+4YaRZajxoaLScgpWls8jdO9QV190
r78otjT/dSqm4Aggf7oKJ99MtsxXfaJjQhag6tTkMm31+dqXqmfvqzZDR8Ru/q+/1oDTZt3Qgg/t
PIFMdedPY4sCVvQ0mySApLEWqeY/i6Bl6NZ54aMtVmKBV2M3F7hOKv02pSK1pGbH70MhJLvaqffJ
ljUoytHRJaAvugRc75WFwByCcq0dqk8UoVpYwja/W96qVzPFd0gE8zIt9hBFlH+mCNTXJMLZ8IAL
NG1k8VrAJeaT8k5apdnn7D4tynIPuzW52+1uWQD9MCj1xbHMNEQfprZBMnsGRYcU2LNyF2jbloOO
O4jk9aVQRZg2E2rDrgOCZcsT5xThOyq/lm7j6Z7ocucWQVmT9kuB0/kUpe7581wwl7tk6sGydepd
NH8XNh4iumgmHyrOxR0e+yo/JxGPaeVtSgmNuf/UAuZ1YZnOyuEL2WgqReryCLxcl4CovO2FshvU
tDjvIWPX4MWoF5NsLWRYt0k6uKVYITthZXxX04+2C/VWSbIcPPVy2cSoPDmpWTsiH8atqcqp56VU
a4YiPxryDBa+nG4ujZ4JnCx5OL7WEnD3Lb/9qfbuPfPmvxXlWo6YQS3D95aCqBCjCawbxhUughSr
mvgeQ2cFJGjvQo5bnYGiEEkeVH7lNQsWGeXJs/ClqyXTjkLtyo6cz4fguYiVZSGgbNFn1GUNCHlV
fBmWaWbjytixR5OBZV54R0GgK7qtSfjxdSgjUH1M2SrIVDb0TMCjPEP92YliYewjJFM1wKnPMScD
kBEHpBc5pzkuNAUNYNTVPTWEGVKYd97997Y8rChRjWC8N4Ai08fargdKf8nMijsmXDUN6vglkh1x
4SR01DVFHG19yvHN8MkS0MExLRclxD7jbVmjaBphg5ROpslZI//Bc3anDWVYyAUUl1++W/yKVAsp
SmOKN+Fx0/8lJwmPWAt41FZzw2f3rIGugmtH5qyFoOKoRINENxirC565Qq35Z4nh+NpKJXBviX0C
uRTJWS3zpAnxWLz92t/eFTKYltYzdT0n+8hwxvdFm4uSSCRG9C7wLR79uxet0HO/DUYQYQfB5Mo+
iIgEXjbAZuO7P6GqqueT/JpG5hsHe4Ypmz/FM0FwpUecOGIJJNUXpal9xYYuJrwYM2TOI9qbbcgv
4RAUQbX6imD8M0xeVTlFcECs9UrXTRxbq6QPpUcbrA+TMlrLVoOxH/2cfH7QtUmw7WQCnVBSyGuP
dg8bGJXlvWs3K74Vs5i4PbJh52kKCPMBkmSkEtvWeO+xb7mk7ThBNJ/mWLhDl9+bj0NSyQeXOfzc
dHetyY9aP5lsK5/VUlqKn7kCuF5WAqkYPdfqimxTG7FtpD8RLk+ou6QV61fFme1C+gMmm2zJP6P5
2K2Y2C8MT8q79MHQ/Q+EfPE9W6MTUJ2aaaq0o47I3DOt0m4x/L/4AwbW+ATLX0iGrI/A3ZN8kENV
ozEkJsd4F1QEmN2JtCGYdN/eD66fT1mAuabfX+QNfUJVBla4cdaaKl+YTYZPXnraopcAY95wNA4G
japMlK1AmioBMgIOVya51t7RKpjIx/rRRU5RDGgdug/ag6Z5yCnjBcnUq19AJWiR5UIhMImj6tLT
asYjc+Zq+3HFKfKXeW/SszvKSrY85oXCuSgu19M4dQYIZAR7uguDSyRpO661JWhtx4M8OQnDd4Ep
DdL4vMCIceAj+EQBZhoVMzY5frE25ef/lqdo6cKZUi7Hg9fbG7IIE3GC3R7roKH9BKfWzU97P2zG
UlSfb6j6EVB8s23EUaBUVGXtwAm1pXdTiMJaTHvgpuh8I7IdR5DLVELLMbQ4ksRCMlA/F/6owdlX
B0n+tgjYO/ZtkzpVKnkcVrOl/U9xlC4U0d2cKwChBPKEE/H01wIRBCGgmFkZuOwNq3mK1axRd4VX
bg9eXhW1wQDEicoTAzlTClWKBrxRKLhhlOf+n5yiEUxCgHA0HsxccKiJTCsnMaBlMlJoZJmzCeSF
01Lll3O0Ygxj1vpHNFIKYY9PuVTgL906yoxygufVynwvvOmdO9IGdqHntbT5XXwf1hMlgSzINkfn
8/sLBhbPl/s9zoBMxYAfsUQUjL3KzJdrZKBQwdBPNlKRlWaN8ecnA7RZ1IshyX4F8fhRRSkSZPLe
HdV6mDlt2KZ4kB3SZz32VU7hoYyXzFNkvCehrEpL71Ll44QbxPS95ztac4o0RKdPjBK+CP2O8Wkx
4kohibzp94tt7uRLlfvw2nQTTpOSm3XYGVhaG2LIywRM/HFH4jIZF0RLLTom/+ckqGofov5g74PZ
yE18ECsEIv5HYv9YUKy6hixEfHL3heWsP4TomdFAVNGZA1WcSkE/HaF7JWtHTTtuZou2gXXuFcr4
BR9ueN5Nb+P41nj1dVR/Eq6bCyNplEod8a1gmTsHFyIicOOO3ZZY+YsntQYAFdincI5aw+LpElyl
WOK84xj4wECJapfn+rVXuFAUzonsNm1hEkErO+4vn3lpq4evnwnDRqWL3Awm0KsA+cy6v9mbUosm
OUGJYY90Q00PCn2quQkMCFToOc5+NgpjUYbj0cXAW2nxd12TXHwJw8Ls0CMo+KgUMEY6p9d6/bg4
nnftjNf0tqVRKZEPsDktokz9ZgCnLPOZF1RyIZd0FQzzkLBv4U5ICDQrDPBnBu4MJC6mzDNxlhx6
RKJRDGUfdc7cAsHfRXMAN1ID9ndoIELDrqAosVUyM9Jfjs1lsk920pxxNXLkwPiUO4o7MrGhTrFW
XMlAyJtQn7zLi8FbUQx08T9L5GPXx9GjKompbEPyPpBoUbBLh8JJfqS6HH5lbjtXfA3Zktykg9ZL
2MnsV0ngtKmvz69o8a9vGB0DkT+9eGee75yu6vX5qTk5Y8kq2ezETsdQCTyhsFBuCRyPjWbbTcJP
lnYHJYk5lm/IlAdwXVKh/U1PCs/AQ2iOLkwdvE7kAcN5YlvGnAIe/VIldJsv32zOip63sWy91ATv
mu37aP+ojjGOjYG0v9Seg/p4k/WvFYdl3vlAtTfqsiwOmwkcwoVv3ujyb7iOx4AnN49qlIa5Q+H2
CoUkQafKwSfnzYYLVksb5ULGZNgeTtT/XWakKzYmR5Q+lByzkPGrw2dzyI22JJPNqOdvaNalqJoI
HayneIATCIM1/oSyzhxULDaZC2fDN9DdMcBg6T5EjFHVpUDjWPBLj+4C6mNLsEB8CxyvDuhykQ/f
1yTS5RGHbway6bFFth05X9sqS3VahwCYO2ZdSmQajCoujILHsIWAAjhN9RJXgrTOBIAjDF3DORBT
f9DkaoIlbLXnF/e9OkX9Lv4ur2eY4K+R7jbwgpTLsd64CeG06mTOaxGFYreXzeJkkeeSdJZkFLGG
Sywp/oCCJNj/3zrEwKKUJSTYx+2GNWMoyu7uBBskMbPhWeXIsUnjpfVOw2UI57prRCZxuDbqGvJG
RB07KQ+/fQ8wlBaMkqdiUv+AXUq++coV5sAYh4+W+sy6asRlDtmPko8ILd1SNW9ELgdW63va3GuX
n7Yz0xo+YXsiz3EcJFwEdpO70tdJTsNTbULN76nuYXL94mRnCe0HDXywTdxA/csyoBxtBKeJDw2b
RE9Z2XAvNp4jzsCGmuHsqc9OFEI9TTwIN2c119DbbiPd30F+0Dn5H3ZvD/dwOnRl7RHytCx2qEwV
bBxpldDri3NexQN6JInCChFzC+e6xRxCQgNl/9bIu4mUBcPwhvxdRkxnrz5nvrwRjGxYy0wFnpMM
ffi3lzuC+lzzHLAH1tHkQPOHOvPGQQ1SMY/tWj8ORKwZCf9Zs9WZi2o36PC2WSnJQb05iapuDe9+
6yREonHRDY14dBIZ3PcpGBdLZ/x4N9JAclYbsjsBgfQzK9X0NHZekg3T3k5Ym4GUCYXq2y7bN1g6
fOkw2QEz+4rPr1oHr1EVsLW5i66kpJDko5VUBUI+DjqMTr+XF2kFKLO5zub/EnFbKW6/f4lItriX
Ps9WekgTKvCUHcK9hHhqKvj6bnnQTpL36kstnTZ7CBHEbcD0SoYvJ8x9TmpFn8YLehC20uTLKw0s
IQDiDmfjdgo8S7PxhpWPR04+e2OOOeBQHqwnN0umui8zREfIW6H6J4eBSU+Sazk0UYxUlwOkGkRv
pZIgElLTayPFXJwH4/hkXawlvWAGrLP5RhHsvBNuFrmOYF5Vv6KfAwp0krYJ8DCzSXE5rchTJW+L
3CfFF5CgOAzhr7lO/DYy0M7H/urOOcwp5Ogt/e5lhCQmrzJkVPDeKtczd28UIoM4hokNV86KfJ/R
qUrzn7+ADrOUW7UGI0+Szg7zuE9rnhP7FGamKW6unwOxF//sjP8JpHQXVCMIQT1RlZGDdbwGMowS
bSE+GV1T9vnbq6q7IuA+NLK0HHI0sOfiYMF+vCmGigiRMH8TKB5eggrJNC/z563oncVCYWtGrVeR
RzHxXYeGHb3033wzXCo85+i4Moq3jNDKqDpZOVL6b4Qs/BKNUNH9fpuzjJgM5FXhMi45Nq+HDRHA
1reCFDbOve+Ylpilx8xNf1tFHb3KD4zxqgyPuyla0q/pGKUYAfNWEQzIdqv/vexMb/cKNo1EemFL
rXMBCy3k9UZd47CmxBYO78slmTzwroY+NdqzYjADF/llL8+FhD/N/PdXiP+VX/LtoBRg9IzTEVD2
nKFlMMN5ZI+Z/fjZy1+hfJPb8LSlq57sVtp+cb20xNc1TYVq3iBdlz70FwwEUEW/7svtSi+Io5WN
WKW3NyV/l7AFGZJkZ9L9PIajp8K4s1r2U0pjnMeXOOsfbFNIvthxk3CWLGFiaJeqB9OmyP1S9W3d
ApdlRjUv/11HvSOytXB6H9OLKyqBX6N7EbbzJtVKMjSHM49XP/h1O9Nrw3yJdw2E00b3FThihkyP
TC07/4MZh4GWQFHZQMfXQMXNCE6THiUNlHb4sv8fNx44CNKOXi9sRint3o2N5PzbnIWaV8zr50MV
gH3xsz5xZFtpOxLOVUNbiz4dkzRy6yTYlM5jxubOb5UlE8UKsj38YaYYi6ir4Iu0wZMQzO6d/hdT
IqQGQ2eNtoqJ/OdD8UeZxyk+bmG7hm6JvzKDhsnsjk4utYXeUgPh5lgBNIRumCJE08uozaH0yrYF
b3ZPfpooDSqMz6qr4YUtBVZyLTNgtRvmhQk0Ehy5oJb8Ruotp9SgQngzJX+hEL8M5hSBm8IutcRO
UQMDJOEzvyfZyEh35nuPPvVaC0HkrYInC/HLK+n+eUpSLqCU1GU0fHH/+DyGNPXDxXanFyKfHDCr
KnTOsl0Kgq5e0nCbSuHOK5hQEYv8EoHB/VkQz4lpjtRAX7kX/hv0/oNnopRlu93I494OJc2Hn1TO
SrGEhQwFsq1qXrEeVwKYx1ifgInAKauciypwLnWAfh/BDZMCLsG2Qb0pmJW6+yx75zixYNMxojpl
uX5Jw+pMdG5o2oRUQTxsesj4pV3Vs5ZZz0YyhrxIWqKLZWozL4s2z1pzd/6w7Twz+kSloha+9/9M
abEvtOQJE3XeIOQKHM0I6ci48gu6eSx8uDyqn8sv8lpgKRP0njcH4UkYqDincE9wmGAd84TbpuAs
baEIteE9lrVlH9OSMKd6OQ7ANam2E3yIP2hKvo342Gj78GqwPnmgSgXdlUQALR5xnaR6RSk0BVJM
oPSVrRFTxY+nAc7eoIyDUNNB+dHPSC7g8Jh2pxgAzesJyJ6h6b+7PdKkfwipiWONooEh+Rqcu9xw
S/6PMgLWbzKCAC1pkc+jsSUGYnDuwRza8Xvf9Gy/qFtEE3qIZ0YrEwy1pNQxTd7mYdg2BLd5UqIN
wuDUnwjDApuexlufi8BULZx/yvGVmMT5Hqwz1vjVCusCz36T06LdaubB+ZNdMgsIKF2xeKP5cOJn
fxEz9Z1c2mOhSnkpt1E8VSA+hyeoHVwD+NCxhk1d8nRv44CRwHeD18kha4NmulcQoj01KBqk/qR8
492vQD2nZ8Dd+MaZBQKfPVxEtISp7WglmJZzz7Ii9frbM7TIO/NjKGOJPVilShHnrqq63NixnpvJ
mRzTv66MFcMNYb4JnEfvUsmjT+o/r2/ZVUY0kI75xGlvTYaOfvERER7fnshiHSAMpSd3leDrYmRT
dNMgpCAiibhV3naGt3VPel2rmJUhOA99vUMWpCiq1MdA15Goc143VOnaDJtahaudp34AGel7cmnr
1OxncrJbFhJqS1oOWQNR2LmpN2nUXTKUMiQwu6IipZy9f6acIqU7JqH81H2VNZDiBHonnx2LOE2F
uRk71o+g3j2gpLuG7HSrXKJXES01NBSsdFxT8Wpyy0AjGT6b8mC3+ToEES/ymrSAlxKjcyxQYcW1
szQ9NHY38ZmDA9LwBsk+jrMh2BNJrA4J983l3YmNk9DWARG8o21z2m5k7NCeg6Fg++3NH30bWrMq
cQTzZd2dbOBBMMX/fR+x2hPShk5OL4bCqfOVoInXP22E47/Arh3/hIO41c36HggTpKQBZ7EvzzOi
NfEiurXSZt0tm3PrOVZQXQXozQKY2161E3qrfG6Zer0Az3USr4AkFs6zGQitY231+uIPBamaJbzK
BX/NgCZ62uXM8y1R/8TaauwcqN76M01E2bmKHSWS+CLtzCJsC5FhN18ZhWr500AOY4d3lOohWN1T
6oN7LRhjhHPMQ5jV0ndBvqPONFV7BMWXJh8TNbdjnkqIp7xjDgbUqZoRG2rz1NO1WM5j3Qk1OqIi
ISKWPBgrZVJwW45zxyoGDMiyRGQtEhP7gY9iRTsYNVTV9QFTBwApDoUZfqtbKJXjkR76Ta/QVhLD
HTPSbg/Qs9028Y3Iohbf4dTnbBWUN3gVPGQSNBdvVgHOTtf19CofcX0hSLgxWtUfOa6oAIvHSxlZ
fGNPv9XNMqh0oZYimSquP35QUL5sw4rzhCOY+vZxATunaEcVvUiXIR0g+SqLrNrwKAxQVOhf13wz
nRbAaMdFkwx8CRP9u3H0HvMFApe734eZBTD8WQ2tv1jV1VXGOUKQU99Q/QrCMJqH09jdWGbvxJOh
GSklf05XYVEZTqOSStDistFUTpurKwSFKi+YeMQYc1fAnEJKfogqLvf2uEz1wwh91SoPZG7m/dru
8tq4ASRKxC+m7P661P0S8FnxnsBYJx7Z52FytfPy6TUzoFORBYDTEfBdiYwjY0tFxXrVgDk/T2Cf
un2SfavSoCoCsWVEIlymoANxFIJHD6IOJQOc2Vp8FOxUA2XvleYFtD/SvVO1ojFE/U3VrfhpxhtS
aVHsV0OHzvm+gdWuVo0KUg55GhJhIaYLuwsnasLEEeodX2ZN0G1UCXo47qFeceFvuAy1TithE7jV
BbITn5do4NBcUu3QX4c60X1u3cIkBYfzt0RjBPKdbgTCWtU5Rb8DBRm2MhfNru+6Xn/DoVj9Keab
PLIzyABkk3D6ippnPuzl1/weaW06tuhLVoOSF9qLeExN4oJLSt85sE3V6ot2rM8JIWYJumhGYrw5
y1cINYhHC8j7juWGWYj2QuFQpipVVpe2vxzm+2BuV04yS7V/C5S4kFcvRcmWV0ubOsgdfd/v+eHq
dTLMra9jswSpI9a2P1OwprJHYYWkFBBQORCOTjkuZpNwz4kw4L2C+qtDeAme8l4uH1Ga8s61Hi2Y
WgoUYN24KzbXieF7itl5jUFUz7RKkJ3bYiSSSn5EgGyJx+QXCAeVEnsiyzXlfwBwPLr057jnQdYg
TIM7crNZlZma0i7Kju0rkjaZw4ufPbZfyfeQKGpB8AZeQoDmpVgum86SZ4nH1JZ/j5nQZ0Iyy5nA
TR6w7JlUEqtUGNoPrItMdeASTGkHAvIGu7Vw49+8aH+L2oqcqiKZuHu1rqGLn3ZlKzalcGui3yN5
9gDLZxu1pv0T3SaILoLnI0WbGls33ur8zd2i3Ha/kW04tc1QSZwtNKQVMv/Iv6SUI1gZLAviV/AJ
HLm5u6J/ditOshIXqEHYEeo5KwThk1yq0BPjlfo2Zv83FPgUpaflgaeKZDFe0Jis6h0EMry4jcpR
FvjLdWWbuVE8E5hufjWV3zci6j4YOXwmcpOupDZpFp58xltQDNibBHDL7yrxpEt+ixu2ExFOpnX3
6NgMICPyNOiKj8oNhAl8a9dVy5dOY7LTUzAVy4ozWzbCGEArRPE5V6aYse0Di4VQd5T6x+yE93je
hgwvsWeXw7gNcMGXvH53WV19x+iKYuzzdqX0bgrbijG2p7VJKcutd28bwdS7I3+7vl5bxnEJXewR
5V2sd4MFFoqyKHhI/mO0IDsFYoFfZzn4sPQTNykbsprh44jEREd0I+ZXfG3z6ZgsoNqY2wPPKmYZ
gR9Fr1qNHx01GSrNSDc6V4CE4iIr/h285Ilr3eV6lRG4Kc8b7ZoE8h7PDqq5d+mlZT3QGpJupTLh
Fhx0ZjX2QftNGbDC2H5uqyr+tQkHe2/zQ0A+b+bmO7LX6mBQtL35BxqmMdw1tk78hPolYapXfXBM
dfM4RYwF218Ip7njYBLlYmiSEHC+PNskRWAnTAa2PLs0twd/h/oWTIz3bBTfcFYIYe7R5hv8YcBV
2fuqRh6Hes7rYmykRmTUMVRitFgD/RDj4KgLRqZbUWRnDNcuJ1P4ErsMA7K5mWIx02JQTk9vUWf4
DaV3/ZuZLJeXI25HROPX5Tgs485a5nmsxTdbWibR+7R+izEl4R7CmJkjvCWNFDf1bCSf3JymRgW7
oMbpOfAVUrzo4pYFdRbOsBVxfNExjBHuegco8oeYuBt3/8bS31n+l3KuacxJlk4jy1G91BQVkWk7
FXLwtGuSJLLzEkyKX6tajxPL2gbskPmTa3jQLjc4H7TUOE3t7ENha/rV0vkmERVUPBeQJDbj/cb9
WKZGBdJJEYNN0Olrti+uSlNP4lDvVlKfSO0G59jcgt59lRwOCojkBN9J6LpOujQ/aF5kEasrYcxq
W+yn+MKRfUDrhKMhVsIS0xxK/oC0vHNdrQErUNgm7+w1MjUd4PuGdsJpULk/zMAw+J8sUCpZpQLJ
0WgzvIVecGhCFFzJJ5p76VFjHGk9XupCH3iCoXhLDRTT6FbDNjHw1KGLUsa/I05atAA+CjlTYYgX
XQRC5VtEzmGszTB6mEU/UERPawok0aVNw7m+jzIxm/MrhCghCAuDNl3ffMtPltDucfZ0RpvsjZev
vsMvxKySeY/0zyP2S1tmpeRZ4gblwjHlOvJ68/Kz2CBwPY4zcFR+ah0uhAo+NB8T+F5tpHqv6vF7
AWBgFZ3yZtSwXRDxZkEffQm2ZNkecs9oAq64xuR0LJTkxC2pSABLxHuU742LCGdCfpto5Q+NYVIz
4s2Y0UCzIKWrclKttXNnoE+HZMfFHFOtWUH1VBRVfs1gUcyolcs2D9+A/8+IRDW+tP3akq95UNex
aYLjIUWXAYameYQ04kCt0j8/zEDB5BSFU3QxiZBEFEthPT+7Gk/UnG9MPCQzakIP9fWmaFf7bOVz
gEPFPLnr4w8ECdL5vcunAp6DljPkYtNFwqk3Gh4bUSmHsSB33DjPrMqIAMu1Rrg2Im3Nezacp3k9
BSYFIIsBiS7Xf76Q9/t2jlmEg7/yXJCTUhDNy0X3SO9pVt826jsjK8wN2OdrXiU53+g7UK3pzltg
fUq3nr2HBhL8SLH70IKdh8JQqQY6wr+mnU0kBGGqy3kC4Zg7PfdkhYW6OfqNsn0mrsAx+zcUpOpb
lKna+S7xNKcDkKCGImTu4IeNopYDHql+sIIclf0XhIEtM0vWHmhI0MutoRh06L73BJI0Es4iQhJi
iZRndT+CeqZwUhdI/1BeI2vhEDkiQwuG7/fT6+hb4W9fbA36Y9e2bLEwUGeyblO5KXa/7Pq0QVip
TS88DYFtCPfbL0Cy8qEqayUL9U22JwgjfNstBb4/vAklUrC/du8p2yizGhrhV14/kn+Eho7Q/0fK
jGgS03oUboa45x+7AATpavIcjje+4X2Z8A3+TWJFKBNSEQIRy86QuzZw/UY8amcqILPNSz+q5z1I
Xy14KcNFRur6S4pHlNF16sn1vBeaSw4LCG7cPXN4uHWWPEHpP8qooPlbds98cv0BCpVJXUDEHtvc
+tVGcLL1YOMt5g127kiQXZ/fWMKvhv1jD1BrYMG+WXTCgbgn1sgJdql9cwbJUIMqfiSjQtAqaQ+e
Or0UHsaiMG2vUDYS2hiOY4fxRR641SDZqY9JW+uzDsfL1CpX8tqpCYeFQKl5q53mU4KYgF8SU1OF
YTnkOgbGID8YSn1J0sr/YFs43UTN30hbGvouXlWUG5PZi3AfpC15Ct8UFMgbgB4a3+I7YMp571xx
0AbYenHeYNHn6NQusW8r4sbGvJSgOwbkV56osALsmhAEjhjubqqAbvS1V/OIzMBtvYv12KAlNM8t
F9Z3ud1NXiMX07k3Ofp8qoGoWo5qePwhT8ZI7SUtjaHYSt4Fw59EJDcLp0cU3okmXxnblYy9Txu9
p+Cp4pKXBqoqVbcz5LVc/Gtg3KpBwKnLaSG6El3oyOGxsixC1riJT4AGgtExMfEGNMJh3b0sLc4N
tak3zTtMjRsAPgCYVVFOm8vNGvhinON1hFshNSs38Z5FpYC+YRnuWAEsZ2KOnLnTEP0w/1MQldjc
jLEbf1ssOzidIgP5TCxwqspgF5ECOkuI6OSjV+ZYO1pMf8TRndv+LtEvXJWTCjIiiZ2r7/TvIRyx
XwUFOeOKg6ZOemmWukxF10bdBdRzYubJ9EpMCwoRsC4G8/xW8FJoqLhsBdpnTwfP/lL/idzBUNvm
nbd/pQppUVBL6R7RAl5khdhiZH4VVIM8bjdQjOXJRhmHLKkA2vIJAf4yJX2TC33N3JxxhmeUIIIL
UM1MfGATOx8yOueavRneesmbA4kjltsqxd6ileUSLCudrDU77YIQt+cTxXjMoHaRk0yxMPF/SH6C
1sZA+RHMM2tv0to5mApWVATASHZIP+V/zkHhJr5g8wWOZWlQ8gR0nfQD9DSZ2VsuPgaCc8ldo5hW
8D8NyZC+DOgO1uc1WsG58ziqB21hUUbMM1LiNlLaQl4k1vWwNLF7Kq5BfLY4sQPRWE8CVpmIRj55
i/6Q2KAtn5TsxQGy7AzQ8gpgMvIYo9P1Sdj8kEQKeU/UswILT6UaqsO2XW8nSvT7+ZN9u8j996nl
09uNi/DwTlvaDEsD947SPxhwLwJsNZzFQjRxKLYsZOxpu1dM9P8N2mrfpfDwI2chu4KG0D6GHn27
a2iGG5tNC51K+Exq+XgMrQH6fElmWX84UMQfUHowUO/tIpYnwPtFx3bduFegevDIa2VX5z19wxZ7
NPSYiU8C6aUHLyGK546oMiCVlCYwy0PkwmA47FHXfUS2i4XwKTOviXgY4Cel4dqjtEyPw/x4aJxo
Fv5vYwB9+atAhZuJlhkse3Za+ezVt5cjtXPHVushLj8DGivvIScyj0cCu0pM6aaAS5O5k5LIyWxF
UEjaB9W7fXoVNqswfLv5kMQwubZ83Ex6p0FlFcmrdGub/sfO3st+k9lq97dpEsliTO5nuKN9ZdN3
wkQuT7tLysKwMc+jG6y6xiCWKA1IMpmWslRIp3cplNrlCxwIP6CKXk+GpJn6fn2A4PRhcYxzyjOs
zN0kehB/+OA2LjNeGN+QrvTfgyMMX7nDgMXFXMukHX4Moexwzb6ioe2XOH9In9HuTizvl4h3W4KN
3u8Caw6o/EsU4UIjpfC48Bxvb4QAAE7dhCkbKPLhuZg9BZpgWOkKg1GeA+AwL678xk0+9msiND3/
1qSnKgSs6RsNBn0aONbfIN/oAYG1luVMrBByWR64A//ffdRPDARjjY+ACwf/7NkNlfa6lbgYl9zY
KIMvZn/80bZbEhceFaDb3qY5eRZQw9SycXobB2Y0oTlRmG/CMrPEJAAabntpTYR8lh6/r2Qw2dqN
7okX79SR0c5/5TRJKw+iprUpLrZ2HyecJlgjZ8cEgQtXkPq8ot2s8ihMYaxyt9lbS68V5NqxRLlt
PmoOvf+wB6gEYro2wQK+Pf+dGYAcTRsyJX5o6QQe3fDSOgQ7mElNvThRBsjzW6wjCI9wxzWnMb4j
VUC0eUFwZUnS6RLhoCBD/zVgWdUih+nYMLoe5Sdz30wxwfx2NfCFbXynIu5dNZ7p1TEJ2x6VlXjc
VcDWT1yJp1xZZsUNBt9Ha9ZTpbiF+4Oq2YixCkRn0F2shl0Y9U8kYRU92b75rydi+6SR1hUYcAXC
opaxC0E+wl5DYDsMwee8O+2lVsJixpan6UH0xdOJWyFxGpNOnDudERlamGjuCKgLQAsztm5fHbaB
NTjUprQzPWVvwZC9QocmadEWTUHMAcvht/U370khKbKquhJSVxcRC4+dxMWtEcGA3BadtTSs2c1f
jdsrPYyW/CWhT43C59x4dOuVr0+smgXvJpO46gr6IGjzcTMd+HlL958E4sz73a1+gfwRY7501vaj
/cmw3fY8g07yoq9M4jOI+OsBsRPp9nCfmpO2NVpIa+c/TZy0H38oMCqEWuAb6hMZOL6Gol22BnKo
ehILDGN8Lbb4ZhQWhHJtg5y1Zby8gx49D+NTZJD5W8sfpw63nkVr417H5+L4yWbUyINcuZ+Ru6cb
Yi9DiNLsdQW6O2/qz/mXahXJkgvfabOAcvAV5XI+vexVvm1A+iw0I0H6Lm7AZxD4kNB9Y8v1JUgG
+rLQPfJwTYReVIx6MldqiDhNWtWrTq7SjAtVaVHzfPf66bPFCEu3E7j3UrrmcEyXznQyLxFmbvMQ
nnMl6KZ7t018vtIbVz7tlOEPQdBeNNG3CWBlVg9T9POinWv4MAD03lZDccvKs51JvpqeyH+bmEk6
hg0Z9HTumr0ynFwx9mD54brKno6rVItdoLLyR0okdvc1E4xQ+aSpHTTg5yuxKIQg9yvQO4Xl8pRq
4XxL/xJQ6OiMmIVgJXhV+EVxn6xJnZPFsTdIgpb4Ci53czNJ01kwyX3Q20NBdI5p1msuZNz9StSI
VT9ntwYE75RKl4brdfdIT9QpMDwALMeMk2cXI2HaKSn+73Nb1AhXMsGy3vNDLClDMuH7ZDL5WHqi
oBen9MS9llG9oZHGnw2ughx81ja7uju09x+ZJbV9CjbQHVC9Oc0FFSVUf76Mw/72nAqzMsxoe6D7
fAR/Im3e/4qomD4aBLZ2thYEJ8VuK1JgvN2aEA1CMY1SNU8l9hggNX1HQ4Y65s7LrgAGeGPftORp
zx0iSywWXR2Ppv7TrlgnesAxhZRYswXCO/OfLbBjF4r5h6sNSo1jzaxLl0SN8WcrzEWnTIV4Ah/4
Mih2hW5WLnoQDNwx1XoPHpdGkYAwCoZd+mULnvhwvI5s7IQbaJpwOSX+L6PZwMbM93gKfjrQ+PAN
h5zQdzb/CUjuJGSGRvX1iyRa19Vegd9htRnlxLBgTsTHobhglvTpuJCyM7kUw+zNwvy4y2RgvUY0
WjCM6JVWpTGwm/RBfRIwA574j3TELoZ5q1zaxedQzDTadqcBeJ2Ht/bICc3O9j8THHH/T2D6Yr8Q
oUnFpFiwDzS/X+FMRYgM5W059FwoRdSK3mge2pfy+CbWiu0Cfr4YRRviMoVhq7U/y2bN+iMh8/Vr
nq1toc9EvQ/aaYznihb+gz44a3Q1CArK8vRUzpxXZMZjCPLFKDquo76NFH6utICt7BxH3a5cXxDM
69yoh2GlZK1mY1OL/EuZ474YhWpYdvbIFp2+ADnP2/ZZ9Z427vH2igGUst1P03l5ugkT6Zv4bbs2
1142ZXBXZgNLYNWVg9sRjwin3p0mqcR1aWci976gBEbxay8f4FTFsCchZ7PAAJze98QHQJyo8W2u
AP/XIdum03sMmvDtlhe2RBVsXeX/8AtMNaEcvmyIMgV/iuysTAaWTkIIV2bfuEK/MRBocDk0F56i
MKvX/UlMPYyCe6upm5N4y4csSFd3WQRyMq7GFBe57WU7mQjhxoITgLLkT5WjvoVXcsB0GIHuoCQR
SO0PnSIhn2KqEQjShgOF0DoJQA/afsLhodnAPkrwIhm1ihDgV45MyBOf2tYyjhfbjKGPbx390fAH
njg7YhXpfHxD9vsOHWZOcNDp6Aoz26e/DvVUrByPBCgytbbCdNK8aYXRN7kD+OGTUe5f/FZJx/hQ
a4995zu39vFOjbPYqCplok9wp3TDMHlwmOahIYtDuI9+dS5FPRLmbK2rBaRX/LL4NsPEw7Gr04cB
2mRC2+VRXEE8iMuYYSIbGdPHenTYH7Ja7QpFmIqRrbKgaiRt9SFW8E5wPXf04JsKLh5RSoS7z2I8
PyBB8CpboKSdxwtOI7n7OVcm/t+vVJkF0Rg5fqe7rwSvnesA9k7QxJGsK/XTwiCqbxhRNOIEnKUk
HI4Dd8Xl3TnpbEsXbcqcSN+MQZrnH6Ng4ncKty5u9+/+6UTHOqCBgK8mME00/inDzSR6jWBVI9b7
cnPOMMG4KfgXije05nYbwIxg0E1u8UV1CPCshDs+p9K16BQMVyBEF8LqJHdkG9F/Tp9fdwYqqafX
9ypA6HvBH+9ZMpcGXB/VAp0SqNsC43K3Fwn3oZoUF/BKlzdqRWjoUnRWf35NO3ROoL1tEDBJvkjE
KySSk1E0PSRhajHWarVxVUe92o2IhmXo5b7P2lob3s2tS2VFNqxwZCL9CfLSzwMY1pv+pDfY3dmO
m1BsZF8ykWiCoO7wyv7qNA0tMP3+zwPf3vneneO/7/Jtbrp3lYW2zfV4L+48MgUIGk6gCFfctok9
9qQXCZt+NcQg3Gzu9lQ/JfGBXqlir22kq00/pV8RbMDOuGNSdUvSL9r38etYeMxGzajSe8W1TFrB
kz93bpqYs9kf5r3A8mmld6QDnTVBL+wkzkXMd0zzmN4LYM9yaf2BgS05Yoj8PPehh/7o53Fq7OYr
gYPNdOsX7l1/n4SeMPsB0DYedWouf1Vsz1KKun9oaXC5P3dEJsbi0JuWE4FGndEASoNUU4aMRqAb
OYEGrmpb6dnd9gxeaFNpNAtBh6DQUwpcCmhB8adCjvdkdwzTCkt3OXrUQ4bdUAg5ooGVoGILj6CG
Mp6q5XsXXLITh6EnQom81+qnYtseraMcq+d7roXj63Lw+xU5SMGlDa20mpPScY2XkpsiDrdF1fKl
VkS2qkroWNCUYdeX1rxR3nuFao32ysEOHjXvKd2XLXLtVKCyjZHnlj+iPVdrhpEu/WsQisLUBXYg
SLRAESypMu+CIYO/hvk8VreLwsL4+gEHslpsqSCoAFb5sis0I+quo/zPFX7AOO0KqIcKI9+CnEi9
MUU9c4Qcduqe5wjVEJxiHZfWoXdqPm0xsjHUiIqW+l3vZkFzsgmEDYGEVCnow6Snurhx+cZkcbzx
N7KdussQ1bS6VMFHx9VBUxfKCLDQhlTB7VH/Cu09wFs+dC/dCqxLpy8R8DwYvmk31ZGCBawp2ZbQ
7GyOvkr3r7UQZBXvKPdAUwRjBszjGqTl3vByA4WG+pf/blGWyD5tr9xoxJQzo6BFS/OPDtb2Y/Z7
R1NaBB7FeVupXRWiFq1KdSgsZZVdKIxB6aa6lEsHLCL0hnRj9Fv+gIVJP1vqw6iykyb4uGVVmQeR
6E0aC+5LVVd0va6dn0YtSCVrIKt3HH+uZiDd8ROMI8OO/p6wSCUXyCEbIL3JGgu5FsR84JMk4yKR
8dlqMVWoqCdAKepQd27bKwjVE++liFCpVuhvK9GtJt7qVpY2ItzNsrGq+2fWjee9qdhpyD3x1VU8
VFcUlFRssZOtBqesJpjV4/hxf4/mtUjdiUZmEOsTfUvn7Iy/iB8asufov5ZMNQZcG4XxvsFAsPGt
oWRgtY7nLf1iFj+FWWH+326ilEHbFViiSeqtB9rkTjqe5bYYqm7TK2Ie0I8vRNYldVT5OwQNuGUm
Dm4UdhCww9rkhYZVOMRi0jOnxIX37JdaQTtDM9oh9YkcGWIfdz2KguPmgENghvruBQs3q6VlF5RH
TszqZyNc0fYEwD4ySA9pm2FyZz+2i+DqQPb2rd7nvI12DUgnDh5q/4WoVpkHG1XCAalWU8byh1fp
vcmbvQOGCCT3j5aZlKwGF8P517sQt6+AW+MZy6PxqCBFFgpTSyBMLatRxOiSLVU0DG9vz5vknAVi
q69roG87a1CnUWW0fE7DUZQXkphriugZrXrqR5NVJ2QvcI7A5lvG5EMxk7YyPAcH/PqIx1BLUI9v
1sT+DqmmmD/P13Dqp1h5LN/I5CuAIrvJaQ2CSTqrf8dkYbToRh5OF+W4BShSQXvr3adrBZktLooT
m2ub6jU01EXsabK9+lmZZv1bOR0O2mz6+UoIYOnJYuPyick0D+lAjmYuLxFPBUWIwu5dzHlfBH1R
bned+OGOKMr8v4VFnWomGiSNL8yfJhKCTZwZKuiI7m7LSbmRo/LS9uDGazQaMWapchXK+LadgEQY
Un99lIeZRNo6kcMsvy1MZpQmZx9pDs4KeCmt7CpOyax0UTZaCuJ2M3MwyogpwPNcCmvx2V8PBs44
8bXHF3143V1cRQCnILjYkreLnCU2xQ6xS2r+6/obQ5TGeBMFJuwq4e2Rej6sEWbta/0tTt30RBAi
t4vZuH5/S5inQKkZoQ/wFd7P6dhUXscNDL/tlDaXHEuzyurMn0z7PD80oDoZH7kpHsRqIDcmKFVh
xroL6DA/R71j2pJWpu/Gk1nnGqFUICVgfR/Xai0jtcw0w3AfHaP65Q5eZrcctgFelQnZVlMkWIOf
9QzgxcBcPKmJ1f8zBpxunKVzwNaVvS3w7yMr5msj70y7PGn+xmjnFvsXuLaXN0YAlVpXkdZq1Sek
Bvc8pvVEwT7ahwXjvSFdXbjixXJsVLSH1AX7nRkN6kUjwnId4R0w0ef3Blxx12/8C+yJRGa6zYE7
FghF3uNYk7BH0w4HmroB21ZUnLKS9w33sgF/IpWXDQlVOmGU3H5mruw6sA9dZHQcsarJs1BN6eBX
8xhfeclOrQ0P/GfqdXpo/IWerAa+XPBVX36r+7nw72uniAKHs2qF6C58JMwHVmy69BybTE8QfPTB
d/JCCBceC4Hlu+AOcs51fXOXpOwBURpZVCsptRzHy+CbRPXl07I9rMDqlFHTVRC8FgiK1l2ZbgVK
lkoa2CIyMVJPaBvqPCH4kBn3dnF6GRDLtkwCqcSZHZFQEXLVa8EvF0OP2ozlEO6TKmWwAAmK21LL
heMYLVIhb3gtm03F35GoEiugJljvnBawwa7iSUZeOzpa32F+AcgSg549v+PePuysvDEh11TCZfdv
eJJQA0woqGtIkfixBi9QEWqZRMYxKCdSUFg7dgv53P5u5kvxhPGmMeULOtlJ/G1ddzO9GV4l4SbK
1xFdV6+re810wyQ5MOfX/9Y0tgotlHVb9coPtQLZiBwvVGeZ00Yqv+1EczVdsi9KXLskz3uPmxgg
XFIyObC3EssRb0KWCMv7rDqC8IxxLFvomJQu+g3cU8dJSjVNusqffmj1vaqSTlKqxPJOIEnPDor9
t6G6xPtnxP9dW1lUHhWd8KatG36za+9TDPu74J2ps90UGxcCR3P0x62pwQOUAF53F76+oyKPfGla
GUlylrTnBGajNrExnigb3ZSjcqpkj/hjVtF7zcDtEgGtxH4XTCuYwW5lOTPvgXTKTyMXTUm/uT+7
dhcj+FwqCjk+eMgNLxMQV99AVsS+Ntjl8WFBTkS4oIRzDJWdKVAYhZdRH9lRMVa24fEGWRpR8+XZ
tTF+toFeoWVYXw5FWT/Owog8AKQdS20asNiLAsWuq8rczhsmFbFJzw4+nEkvxwWk9DOvmKBMGMqF
OaKgP9KifpHg7CiRzKJVwgaGLCQYHciHc4+oZE90dggVakAqOI6GVjhxzgUg9AA7HnvpNI9i2QJ3
qLE3sUdox7Qf8MI8eJgdIFiP7FHE1HkwAcmUdf+TqIpL+O4vftW5ky/mXfPn/et3FJxnw06+N542
DhU8Ov335yHQaJ5ja/DH/gVv4yjeznPMGVF+NU2jqAhfgv63HYNz0RuIlWGINp8wV6+qV7y/b/tM
Bm7E8WW6VF94uqITHQuCmObym1jeEGe/+78ui2wvJXZetlA0zKG9iK6g5yR8M2vvy/cBfQjrTzrd
hg0xiUok4nlekuB9XI5gAU6Ui84iKBzW3Vz0wDU9AUCgcfdBO9WYPMY19r7oastii/Zn8PgH+/qy
w1RKMOV8gPhfhMS9YTf6sTeJo30oD08q+S3P9qWrpvW4wOIwxoPg2UmfKtQmWY2Pr6jaQPGadNVh
0/mzH05JRvUwpksAT4mBeg/wpUVsmcfE3G33fYesrwDRrDSedBLUtLQDLKas53s0NdzCsISs6Ahg
RxIdtDOAS6qHuTHh/wsIVtFm9RInaE2uK9gpG5v7HzaSWx/xNkM9uS6NGdUYq4dfMFaLitYTFWW3
GYSCGAJTCD7/PKOX0HTcb4WqJAsJxBbiM0hBhDyntMVPD3s0Bc7hD1q6NjxKLGVRvMcFj8+S3oE2
KZdWn1vKdHB3NbR1aJO0l8ebIKOmw+5p7ooKWJHfnF4Xtyvs09KujnTyumPU5LWVu8Nf0n1sdA0q
5imHyHeq/gdvOm3AmxnvfL25eZBhnVz470k8e+Vedy/EcQtFHID+uk3DZysTfUPy64O0Io7VGuJ3
rklfgISJ9mikl1TI+jXpo1//u/y4WhQ0hGlbgaFDEUUR9nwGvtp2+gkvDSZiBiC0DJxfdm9oguGd
sOIoJkg1p6DLrvewNvLQnRij+A6IHQRul2tLHppGaZKL9OLOgJ6nWPtN8IQyzL8a5W8qffUokzcD
gmtlr3lVTt0/g6O75j0adkUdgCchaF5RwplM+uEXvqVjjBsLKlPDyGTFHDf1mm4d2w/8dvMIT53H
OfLpxL2qegkAcg8aIMfMvkQRc7nnqB8Wjg7oEdZsou8db8ZYZ0oQRV/yYUkZJ2DEkJmotjhrzoj5
IEwrK6A/QZs1JbypTqIM/lHaJE8wwy8WD6uEsca3rWCMXU3mC12A4wlwfHIqeOGg74RK+PlqLfQJ
lv31/cXKHs8bVv/3SVZynL21atlBhqNe0K6X+BMxZSba9+un07QR+UUaxsff7ro4eBBcnl1GuP5V
3oiTvTyWcAJtpIiy4ro76srUWLD3g+oOmp1oY3f8DwJQiFMATQFrE6+HC8+dxNwXYFRpffMxC17M
deOD94ZwWqIZRpiNO034yat5Z0XbhCBa1tdm7yd5yHWaqIBd1JJ/RNeXoCRnKTVDPVgJOB6rlN/1
K+3JnN602XqqMeH2yqt3M/Dm3T7o9Pqgie/PkalFg3bhGasDX+bhJ2jl3G107j8Bed+squW5VssU
2hv840T2UIbgb/yjGN7Q9YyFQqbbLDbDDUzuC+LdSZl0aAv8al21Mbl3xNg88dXk1ucuhkPORJRl
UeHcEl65yG71zyRp51M34AYj7UUMz1j2EFJx4GWrcRvEHgezArkjdoTjM3pd36jEGgU1DVgeuZD4
3WPutmKZCHeX1ghUfKNndUJM2kXMmUzQuGuNISHIVLF3BWnGziLEQo9fY+h5F6cPg3R9Dcs+0/dy
RJ91WQGdXFZ7oLvE/+ILPh2cNvD7W1VsDWksj0Mv4rPKisvivIRqD1bF5+vs+8+O0XPBwvfxgIZa
iFS23WH4/xU88bH1VCX5I4i4jq6ZE0HfRwm7CP+qnluU8SPbYIqUORSBZt5RJ6bbKS3tQ9FZOflE
xcPeQJa0kOVpvEH6n9n3Mba2U7xDJJj/XOGcLW3esYnCwZFzz4aG9xPCpEUiT2QTcY7ykMubiog4
64M320YvWTC4vq4nfZvkn7UrT4aQhvGIVirqUd7FEH4oIg4LYrBqF8mewZ+ZDyfB/zgyOFbd6gP/
ypgSOLr0D+IN87tkvkqnodlD6iFgH9H81UQm1UexCLuYG3QhObSgG+Q4L3Bg/wEdbeNHRB4l1hQm
rrM3TxanN8qaneHzOMOBDhG3F/cMHeH+6DpT2+WP/ZpSvPdZ8j1EB4aP5zgSV4C3CKV1r02dYI0K
Z4yJDfdaNYVHaMU2+cweG+hXbf+EYxXgIJ821mWMZTwx1ae9d94BhqkzNbXkMuVdl6ApRLPIcGtU
wCEfwp1rR7gQuXSWcz9q/C+ZPj7GIHSoaC+p5eTF7S0o8pRlS2SMMekKvU2qedVQfoJa/ULHjqbf
kp4IUmAYK92CqLLEttQ/JJqkNgds8AdkCvUDY0cXOymlAD3rGkHZjlb1OwUnDk8VWwzQAJlsNZF8
C36S9oYIOCyXR1nvAbgsvOLn3ewm+Q2EX8D3dvplse/B1KQfHmltoqsSHQFWDtN5tLuwl0wAqsP1
QMQj9UHAi+zZtZmJex2f27lGbWMntd1LBKMCvsD1oFbgQkF/NTwE53S3iexGMS0R+989FPBAjR9Z
fv00lXtL6NycO6wAhNYdo39JE2DqUHtiCdxN81yVKIH11ykJloUtB3WNeLGeCUo4cBkyXMIybihL
1WzOhgEHomoyXsj1/Cj+ujs31N4VbQN+JcXTVaGVntEsudGG8SDTNxuzq5I4C/Zc1VsXNuZZVeFq
MTVdHQGs8de3ssoNA9/Cqc4BF59ahzCRfFLC1VEJHgtyLigQUNtsA1E/C2a6Yi8KuYqX28COgxdt
neILBBEeWwVFBQSI/H/c3MEMpmLTniANeILaTwPWjPpnFiLOzAGOl49uz2CBudIBUZXc5RtQAGWv
m5kprLTxx8ajhZLbTgPS6+M2BDPILR9LuIVpu9HWQEoe1oeT0BIWTGBZFopM1HY0wZVSPFBAIdk7
I5V1LMaqMZQv1BhuAro6SfZyu19G8DHL6p7tnrSQOZlc3L+qzV5yOmOOUJf5+gktZN/Jb+tuvuc6
XWr7mbKy7I8H4YCKSdmolzo5/H1pDGBiOQAidh660mJd1IEhqsMC3PmQDMn4LzxoUokwa7gPaCFK
3hugsGFEleQ+23/bNo1BsqpNAfC5hbz/uxKIC86VX7xwweukLhgNiJLVlf+9XK6bxZp8x8tEdtc9
kwpML0pYVzWHZVwBhlnJkNRkxhjFV12jCGSCiGhDXZMSyuoXJnFubgYRvrNex8KjuvMziIOTKGy9
Z+kdEJMGIPI3R8wDok444fXWIqmvDv67r2kBBsRcZbUgEZnr7ARAmYUCzXgs594M5pvs2Omy+Oaj
J/C0gDtb5JRkVZJKTOg80YH8PBOTKzOANkSjd+w7A/1uZsr8oJMoHvqw7IkvOTjljCtCXy3dpiR0
Q68h1VjfldyznqGQoKKjjw6HY5n9nt+arr2YaP/UdmVcpFHdPvy4Biau0z5/neZuT50Kf9dHfUvL
u50nMXkxsmBTgOu389qMu0UeRjqmAMfSnxoXDT9BH1OW/zpXHAn6y/R6B3XeZViphl5CPm06c+uh
j7r8L3qWn7SbNnO2yJZW+Nrm9g26jq9/lEMnn6AiuI3UPvfEEg97ryolxgFKCOChCZDalERqIPsg
OQ2QWZVguJHFquvu/FmaO0ZMBrhjX7Kx4NRTHRnf2ZUBEdxuTz68APsRxxCmhY9qqZ4YwVi3dNlH
ZLCVM9GodXzogs1dZDwo99y4tZ6jlez0Ln2G7uab7Sjqllu3+/JgIESHoHDxBAn6m4ME9AtLXoOl
6+ETyjq7z1h4m9S4bcJ4C9AC5t2hSdaxhVtedmNVTaxpuH56P80JFQ9HdwigwQTUox6SbPqBTe+B
D5Ow41n4Vq4/+h4oCx4AmoJKcBP2O+qubqfcfiFsnscGZoVzge7EVzIrivSF3mf4l/m5tjQMH1Hp
HOGeElZifxBLDcfN02S6v3MlpJdLOzuueNtAjG1grUkPRf88zXZKYXzhoTrk1D5EhaEEdgOsW5/F
LPkXyUF+4La2cjur2mbdNqxQVSHNP2RXUpMP6w6zndo5z+Ps/llbKGGHEEeGAjJ7GEsSXsoNCYEI
C+VBcDPDrq749dmauCGnb3ZHDC2+eHa1ci6fXZ53O/jcD3ebfyN7+EQYFVBvqF2NL6HKC4uqX8mY
UlJhhniu6xH1O3iKD5toypSXCHe6i3JzCxkHqL+Gtf8ItWu2vP9eih1jLFDLjtBzo7j9nJ2Vuei5
2ZPU1WB99z331B5CLTSG3+B8OzUUFJVxk4rFoQ1ZSpJaNx2qVAMB6AYu3OIvbREGGpjhGhPtWDAc
VdIlJ/RfITuEghT/r7dt9+Rz5lj1el5Jp8p6bdxkSqOzhCLHyITOGY9nAnfPIWxzK1B0l4hX6pCg
fHvMPYgPQZqFBLCR/z1a5WRFyC+BZBcr6uks7nowkCs5ISqoF4ubwQx97fzhihzTB5siiCo8BLKp
qZ3dErmmr6IC9y0K+Zo1+dm3jx+ldYJrgQedx64GkfePzfcxadDJ/CJZtkDVo8tSpEXxcImO/kWy
34C64kAnt3Elk7Tza6+sJlIWkbS8W+2C0XDugaPzv/1lC8rG497OKeJOMozjLJsucNA5/rRAoQYh
e7sgepXptvBmHzUUJxVPIivBRhwqFIBcyITOVnOw9FvQ4/Cyaiulht6WtsaQDsJm2aLy5MQ07lH4
mWBv3PJ8N84RCgh/cx5dlr/JvZATsyuhhzqPsmH4eNFb43fvRNQmlPFIr+cIASjaANWWAv60hwL3
1dG2PKmCidBqtdCa9OMyBXVGUMZsJmC6+CNeEdDpzG0x7u5wjHL84h2RZ9xCrl9mR0MPcURBk+o+
5Q/mE48xafrPDoKyj7/MKLuW6Q1utSmvFKjrFxYaYPCvhA0uB67aiWdt5pHATttDHtMS7nvaBk1/
J0DjTVlDr97wkxE3Lsz25k30MVHVJwe0yqeggw94xvHgQcmiDGM3a4U0kH0daOdm3iOaqmx2rk5h
tP8VXEhSazcFxEMJsK2QOPvxOswJgB6UzEvwiCd5nVbrXPjbQuir96vzt7lMsqyVqMHruYdogH3y
8Qb0Xz8vTVq5XBFz78zDCvsEH9KMuYAGRjVFZpAgevu4+szNlQLE04J40o7ZZZg8TwTGZdhzvgKa
RS1Kn7d7Ve8uXd4HrclJWF0WEhECV7JFjisXga9+NgwWCKIphL3FEi9MrdVCFR5U1dLhuRPp191t
J0OKgam4sioPfEkvpCqC7v434gtsMHaHKw/FCoJEZkCu75uqHPKDjw2kgY6ZJ0ReJ+VNba2qLc8D
hfhbjG/9Kug/KU1D/2DqdXnsQSLAc9pyJ3QDvPykdJ6Bcx5ijFv/KI1TeRAheca844FiVlw8fxv/
2rmi3SlvPTEC/Qi+J6o8iu2r8GU7O0tEnsiFNHoPJGNGz32DFj9QnMYY4A+iZNM6XF42ct3RqTjL
B2cGlNkXDn3DxPEs5fgwdL7ZzxDwzQMBVw/8qUtx1cK+T7o8r3Fls3hxrgxE6saevMfXzmLSbjMr
g+3c327BtLo01UG4Z+VgPKtmBH+mHY2U/+O49kg2IjO8vEJ4edIXyG/bkfcEOjIybO6Aw+3Gz4ew
fm5BQ3wIwKOKvLwf8AIkSaJIz5q6XoBRXmk4OcZTRgPSC0NMx4oPHFuKNXC6p8PVfYJta7dxI3db
fesScCvRUWHN+pgUbsM1rf2vbu4/2IJP3ijNzmTHnngXxNkDLr9DoRdwJ3TiRWBuqUNEYjH1iCCx
O6QnNd7HSWg56dWHvdJ/gMzG4ZbFBYn7WFoSAEFsdjl4935vtA2JaoqG6Rwc9d9boFO7YKa+j5U2
/WjFnx7vOGGP8iRG+B1uwzckLGu+le0NoZRh40BTjMxFWiYfgtye8GI6NSqROGrGJNrDRBVmHvK+
8o4xyCIGr4QFTyySE69iiSWoIyeDnycLB+1C/OicNJtW2fVG/NdG3uVFZEC6Gs+pLok/kYp3frW2
+sQD/T2nnBZaYQfFwDVX9cvg7T4Ci1Iw5F6c0dl5NNs5xsccmxWv/KLHi+Hwj3QA5SiBtfWXyjj6
V7WV9efg5fzPBmJDc2aInjnBhGsWK+wI616Ky1DeXG2+WHUdVl5onlTwJBSE3GWwcCx/+zHiQ0tc
DoXfTKhtlUlpIitp5K0TfRcFen37oSXD9VMxk7znBgjXj6SiUjlhAu4Kw8xb+UnaUscGl8booT2D
U37vzlLnQqbUsneV9tC/ptCDmZcMUjh/NRSkbPg8zYVAXwQOeLgAlja2KNhu0cAVWyitI++PeSJz
NTfUaStclUyP9HarHHKtZcfI9x2TFSB0Neb93qJsoT9HTdzdspmGmppiQl4eux0MgLydFShEz4iz
gA306MyfrrsDoIpe9GQShagYTb0ZR8Nrd19+t7VV7GoFf4S5OnMdHXrxLppO/+JELBACiPGBVsw1
PfnpZJY/bD3f7m240MyhHXo5mmdmC1WAe+PhSNDHzotmuLJ7twokgbM0H/qK9j2uMqNO13nRdgAt
v9paBlv3PLW9Rx+oXNlFWSD9SPPo0jZCrQe/WLiBRK7FdgUMb5jEacUial+Iyu8XVY0LsZ4csDAu
43eQ2+dmPfg4m8aEJVuuHeqpD4yLZFsMh4w+haFmNSZTd9W4Gu5NQYCIfeMC0BQrmwGDGdxSqzPW
uubgIiE/KmBpAm9f7OhogGwHrKIiHaon1bpRMDKnMPyNOVScYjj9JhD03qICQ3zvX3BjV2/U5KlH
XJjTwcESwMJs5S+ZTsjmCsElEAfyaZrqulcUaOlRJTsFUTbrRJ+Nm2teNoKyI5O4bhwwzNcQx2Cg
vbF4xwUELPf+xXYGUuk/+jsECZzbc2wiC5X16WVaPJhQH3EcAWjcVfjlCd/HQhQ7CxwVeuMUHDRM
+Gi8B7XKluPkjX+7cdYgMhA0C1ZPVMNRZg4U9ZuKnqQdyKDIGU/3zLQCbLjJ3li5jST4Q8TOWa6w
uVdENjvyf0pa110jTY+DIMuHKiPAbweK6WTIskCwaghc3C7E4VFEEUZiB8sWRYtfrCprwEawwgAC
ZlTXPnnKkX1Vb3TuyxmcyYg0QMuJres+50UFLBopzniiAR+b8j4cvzENbjlwvXK4jlLbhsql3vpF
mklyturJcjjpOLviIDV7LCPCGtQxoLwtvrLj6L36vwOVzXOaikv/2QDlvJILoSWlSgT6z4tEcA+a
ydWwZvnKs84oqkD+J/zjU8piHyHMa2rzTHmvtEC06CTJDDXWDBIRCsZweQJRVA5Vr+A83n1l1Uzw
/gRylN+np4LWi0rydwjzISzIFE5+5bLhtKiejMv1FaUJWMMqmTdM/PLi8VbqLQw8FOJtAZDrVQaL
0RFW+1oon6ijGw6ZzstiX4uS7MSZoz54ynjftXad/CtC/89RKdhYr9S+mfY2bUlMayI902gecHm3
NoVpewqCyAkmL4EckAH3vzzNTHj0N3WFkY0dpjjFkJU+uk1Lt+lbqaASEalhMipBwNRWQDqBWaiq
bnm+MbVLaAUTUT5UapjwOeRYCXibp8xjjHmnZ5k++QYjEC1FTxdW4nmucW1Zh/KjICKWLeBIR43j
35XxJZQz6sl/pnRdlVEr0kPP1+8z1XCW+MkVAt9AzmAaaxTOpuJxHlnXJDoKI41HTDtdByc/wrYf
9gASx5iBT5FE+Sk5eUQJv/IPvzuFFVs9WMEN72gpHEbTY6bUd6FmLqLMbP29rrC1tQHyWa/UcMx3
2fIh6xOBdShvXOHOXwiEcja05CSVy6eZNBtAYe1ZrWKY6vq+Emf0I4Hq5AHtVOueoNLGlnN49Tdr
ka4RTF0hy6ZuiHmivngDsSaochGqQTtJPB17PB1Hm3ClEaNUsDG8TLx9MmALSDaSR2QzSHAfib+x
jiyGy+It+H9iVWlHtI5kQN6AO4t/qCoXxfEb7BjuLkP3IfLWxwBnJrnP5DjMQhrsCp7GbaAYK8SM
WIi5Uhm5K0JZW/Ln3L+4dxaJ2oGiY7pyoB6QvQu9QYiYNQrZqtVd4EQssRwrXY0dvSqzBfCwP1q0
v2OP0Q8ja9Buq1KYEIPmABaBLrNAYBJUmilhN5g/TiZgPlNJ+X+xE6qf0+Dasx5F+NC476IaiJm9
aOlqXiYI9LwJlTfn72/06pBHsFaTeNScNfEdN1U2jFuZwRW1sx/MK5fguN4tybT4PTngO+izbBzp
3PGY5cEeiVOjrpX+JDu96cdr4U54Ho2tyhfR0ByZuDn64qPyPEUBD3F5TaV9juP3FaiAFMWdbpY+
oeAB+wV10LUUgtGNQRzhLJQ6ZpeuVfNTxuFfPmbtCttY+VUD1QGLbBgZeTiXpnMiderViW2boIFd
AljOVASj2qo9Fmeem3zNZvlFpGxlypYIuBk334GLljvEdPiF6XPHH7i0YKUxhcFkiBSj4T01Wz/k
wFBP74CJP6Xfn9OqofWHfOu6sfBvvZxRGLuKw86g21CXB45pdr1HSCxtIzjfSBLiY5WYCMHOZV6X
u6CZkBJgn754C1Vv2J7tI4yiUBKvQFqXWK4AX9HpMratVqt797L8eLbytmSIFgMRaEXuS6zzR5Mf
lTY5vpYiTFPTOva+jA3U7UMB3nXjw7/m1tttBZpPCxWw1AmrQV53iptUQojo13I9dWU6zB/4F5X/
ShiLZbBk6AZWEBKrNBDtJxGZTrI82Rgaz34h4TqKXlfk5PeVi0GgOentWaN52fA2mKhxskiW+YD0
iL18RHT4Lj1I5h94naJLZFxdKqoqVWvx+j/HK2jji9+otKMCAL5EpZMUSo2gnvJI9Xg9arbIe8EB
z3whVHmbBdzZMdxM8xbjnm9cdQqnFfcFLRy4aDA/LZWexZP+jRPl1YoFw/BBZnZFnnD6iXwimf66
/PlxjYKIJakFg4ouKEplhR2bGquvqnkmeH8L1Simml74piTNZ5AdA+iLBQUau/iKtcJBS1/HK8a2
X/qDxdiBJJo7w0ummF1KAe+uKCPDze2EUHUpP3KzaJMv+MsIeCqS99neJRgncs6PNwdnUtyjGyyC
w93m4xRcYG5P1clZxOcjKtM8jchC64aAwAOvozloS429L2sWmEkweeXJIc57UDuIZqLhjqxpdeyQ
SGbaJU3PK0XdOgAxsXiARyoQykf4NPNYF8IOyZchzCKPjKWnlq6e+DEQpeLVBImAfdm2iz3bwJ1N
eLIQaiXXqenZLU8G8m2zXmuKmcx+cZTLNbpwUc9v4nM2n445HBMci68WPKYYMsAjdqTbqqMZIUsW
/gGuupz2hxffq7sHmhKTt1yXf+MUVg5Y2iumepg29qRMvk1v9utaQODClpjkd8plsTlkhQJ04H9X
vQnhZZLp2OkLwa+OHr+tfIAecKrTtFlYqUKHtJog7fILXCd5AEZfiWrXzKWtnDTe09l6KdEBZ1pQ
G1K6V/ioFzj4E32Hee9A0gCwsAofCJw5+rugwgcE0O4+1YH1ghgewX5WrImlIO+MGePxG6N6jfZy
7YSwHtScITkglgL8/IGkfdC9hzHP3fEg/umZtT3QcGiZWQEc0IytQYFME1l+UPIrLUL4T9leBklE
Vnng9DT3fH0/cTCs2hjSf7eOJZ4lzaU6EcMiHigLmPVvExPyW6K9Wo315qwNu2LWwq546rXQeo3M
nHU62AaxzK2pkIMLBDHcbZ2Eah/t3bwpCHs/i0yXO/WSUJYPIpHERwpP3qBnXybuWp9TvjnUfRMP
xG92qpQFzRzCUeFrN4UVxy2sAR7MkwFjmpjuU0aPE4TpykTWayBUDGJCB54php6ACOvwYY/VtfFC
FTSklgIbW59KhZWSTt176XZuBC1s7g5QmPp780h8Kx+g3CeUWZL/BfF/EBHBEBQjulXeU4Va8XR+
PFPuOWKFewz0AUMq2nbh9ui7TrAJnq+rgNAOO5pkxvg1EKE5lfya8e4h1KccJUt7uKkBgiGHYbmR
ylP0vGFQZUgnmwohoXfbFAQqEgafl7M5sRDvBavR+SO45ET46BUDVuwwlnUWnn9esPNcmmr1Ng6y
s6+BMSyVyhYQAX1M8shnqBkIEO13zjzPVk/rUOveIxl078+oenyyM58x0Gd+hlYbtPwpaDfKbm7F
3+ovnQKimdW7afPr/7h0nQWldVsuqSjV6PhPtZ9nKnmc5JuhPbdWtO6SD3AYlq6E5ICah2/nb14p
HFam9//kC0ILd2zL9bZwGFpZhmD7+UdHABTn5qISFQRGGcxg3zZkXrLBGYSmq97apOGEdVo8MXaz
vicH+0q7h8xggs/M9uJgcwHL3vvTbDz9fwBbJ7rJIm09Ux/X470GqsTOdA8ZovVrCpSkaFGgKRIw
GMLMDKajYJU8GGF21BPRCl/LVPQqqsOA0ASHSbzFDsb+jpVUYVRtqCSSFrtpSIdQNF6D22GpZcqr
W08fAGNP3uDAYTQ2L6ey5r+HYF3ntMP/rF+KDKkQ5TABGRainnpUasmK5xxd78ekViwy/9FHDoMf
GGNFSJHluEy1k5D1qb5KE1CLBjTIDQ5t2sFhPpsmM0WYVZJK4f0tuzTGmiAgMoQ3ax8ZGkJNnSNk
XpmV2rL46qbmcXGJRxZmvpFN5sK/mVZaRNNQOk5deuWAulI3/zUmVh9H8sjDLUAoxRZyFP8duY9H
Penbw7GaUF5GlE9DB/ruf4bXC+XwjFB20woIFiJeLwXm65JzWiGaYeGOuAJWmc/mSnnl9xBlAYjK
SmPYyYbXuyllDCMCTJyJInO1Oech9fGiyDGPbVnKC6TGjmlZG4M3qc5L0vfbpaAFPmGgab74Gvyo
PAaH7CnWgFFtxstquLMR5IINIu7DLW3DNoh6neK311Axl5i8ZLqPtNXD4goXM9jhBiELNnlB0kXV
iUqs4RMvb4qtmHYR6600ETbQPYYRDlj0VmhRoJSLzrtjzV7gTuSAU1FcidvvFF6A70PRx8MFupKq
9LGntPgveVJ3ADNatyfBNRHj13EOld9dvtMMp7huW3PAUO45s1A1TnE7ZCtuzRAYNZ4juaTlQUyu
5l4umL8alBnvRFmU4rjfFDSnnR3Xp+MFubrHktPxab/eT5Kle/x0/9LDXT7JyEGufnV9M/mbuppj
h1WRQuoCm0NymiZ/vBWXYI1B2q7RBu1luhKo5asMXwW1Pm9BRa6/3dGqRkl6CkMDy4gaorlaqXg1
0UWW0/wME83cYDp8ZLdFiNVnwcfEzvDSZgfOI4LiunOdnSiZpFg46ScmSIY0b6twNYJUAwX066cW
nTvbZYBxmtDIscFSXkUcTH4mDj6kL0qZx01rR5OiL113G69YkVcU3k3UmN3dm5gW/4T4juVq3raU
c+3SDbHDpkWgxKOwnNjPWl1pgD2LfB9hNgfDANiLVy2jqrfsiiVmF4zKs2npSrFyMvun0kkRQtzB
ZmsrVC+GI+4vYe0nsRjbFA0cYSHnB0+RYga0QJFPsdA2dIHjl9J9gQ5F4IQ6ZkxcFRmBmJhioCOq
vxIC7LNG/1qDHuyNOglFyZiVi+bOGQtiRZ0Rncz6lRpLAdL3N+/NfEgBHj2QCa9NY3KjzuE8kLHD
sxsh8hLtXFvBiILH3jyYn9PlhJV3rUfbduUJxHudeJoZWEqi2ToL+u1KeKROdagEUK88GVmzF8kB
d6HhN8d/KNa/lSM1jGwo2EMPLE4wrBVhIJkqZCtQpkdBkWZrnhG5rA7AlM4GiZo12xWDoZyoQWVc
dJT3vJ4vXts43Eh8hNT7z/ANhrRK3Fy8cGoT9HVhAqgg5PmB++7d0wE+6fIkIp8AclvP6wyIyOlP
e7bjDwirlZ4RgBX6EbgoGFJIkdi7+3H23Zjjt8AKVGEzxnfjUR/eUGgXhJdKucLgSSzn9z0u/g+b
+DsHG6rIjVkLjNKmjpL6x2CYSnwXa8CxzOKuIxqx6o3QlIMTeTx6zmd4leFkMkoDJsYfNmX9QeDQ
4XPuAEY7TEBbzANycdKCkcXf4SD+p0EfhcCEnvj0CAW8uOQ2lJBUVsuLB3dbFXZwAESEwiqa3pzQ
qTtAtOM6DfEXj2XbleUGr2F4VgmryZitVWkXTyMNnaAVkVgwf12wLegqOrcM+yTibMtap4nYekDs
JQWu+Z8EJxkMCWpb6Fjjlt+Wx66IKavPpq41d9a9USkIFM1+0Q/8XOw2AONZunOCaKxTP7p+MQpe
89oOiBDzL9e19i0zR87kYx5MYkslyJVVrlIATPCsylHO8YNoW+IRcRgGrQoT5vfWkxdit0qCFh2A
QHKy4Uk9Z9A0eV4jxxmnEa5kayjA7RMBQ1XI0A8sRN1CCnsDXryjWhCLvu36VJ2W/EQsd/aVx/Yp
fzQ6RYteFSou7f3zS8GPAaGRswwgR0ueUzJUVcwTdNUR/8uV6MFCIkf5da+RQVawFd9HKRBQfUIM
8n1ebhtON/P62xcFmmues4jOVSpxANJfICfD10NbEsD7lb4F99oGHfSupk8Oq46mc/ddyjxch1Yp
pIMWARBjp7gvO5z65kWJsPLIG2Tf2HgCHYo+rOtc9l0OgnRLeVUqKjhqyYuEM34VKWx3j3ox9yI8
2kj9RkVKlz2vtx7XIZ2pWMwGXaMhhKzd7NmKX11k2dH41iVQIp31rYP2+3XxCC5aak+6cJ7Xej9Q
r8414BOdihZJACwi+TnfzkJSsnRgTYGxcbv+YVPOhcgOyrIzffFv8UeGWjkSnpDvn8ZM+NGwvmej
5CrFa2b+Nn6NAmhy5hNqhy+SGARwTXljSPgoOLG5ux6xtxKZqEaOAecmVad6tZcG8xV3sHC9RK5b
qxDTXlSoa0UDeC5B7/ESgYuSuAe3p8A0NjV7W9mc7F79EX6CJGl+xyls+G+NdLK00dcTh07HGtrR
qztNnR07oznmtrFHbqUEk28fktHhpnk89HNm/EmLRhG/FqeH1C3FAQLqYy5sX01oQ24G6ngu61Rx
Zg4jOq8AoSav8C2fq+1WR2vYqsFGIGqX+RauYr7t1YD7Olv24nfS2WrSNEhrPwSPaauJHfMm06vP
PtIYO/l8lczd5HyEseqwxDa6O41vLfXliCM97V34RMzdtWoYopDS0Uvjj3F5CTXFiaO5K8Q5ddvT
0a9WEq2PfuKwO3zZflmJMSL51SQ1XmPebfYsayshI/Vl/hN1ei7jo0cuRr2ogb5J6esB7Slt5Wtw
bWslUujjQAs+93OiuDw/JmIohtrec1BVrvKDUQNwb0JMVu0OMbHgIVAiTkEl0NCi7lqYviHK8Dyq
8BZPrT7Gx9DOwpID1CrHlZqUdD8wnxbMPyU+YzPdZmjBkdp8XQkBFkOTVdo6r2wHi7iFohG1ASAm
6b0p4KWriuxxwUyZ4SwnsFLQYDDApJ/vSCQcLJBar3UvixnCGrrKteuWjRDytPavpIxxEeSsoCd9
gGnrcw4zGSPu8Xrg3LbuyowySWjqNbzCTyv5Kn4ewONDflCjV+p4zpBOXKhMMA1uKYBuaEVvwuKW
Qyj3eT/RcDLscEeHLxYUXjj9WTUsgHQiW6dzaLw4OYng3jvAqQ6gmUSok6v7FgOL/8gB+UEGtV7i
9wvtqT7L+ov6/jsrwLAOjIKZ+Z+B5p1p1UZCrNiqaRiWZI+mARlp+Na6DbnMXLiJJJIZO8ku6+3q
TweniDQSCmMndtkxgHSztnCv2nBXIcWYXYHP4zXCgGIgNAnb8UbaEUU3ESvMgjGT19TOlxZyjizP
rz3RJoYjKnEG1chAQg5o8cKHgQSdzMdFyWsnXHQBiUizykLiTM2fmhJmB8koclTr8faR9nkxczMR
5QA/8HzzAc4pZxdktT5IVGdG67NfMVQTNCPfNt/L+STXDmRB2FoYZQxHeEAtow8krgABtDKmNgzp
OUV+uQHs7woeZX7EQ7hzjp99QhaJ2kQArHUFvolRd591ha6VSalsGnmCXuu9gKBMyRrxbl2ot9jE
IIPlULqduWCBGlt844IH5+tu4OZccFf9o7li8isLUruAXlk6F593Uu4PfJlGejDhtavN1hZ4kYke
3T0Et3Lrm/02r9ct9VsXaKKyzk8QGjV3rr9UUTTd1jPJbaxQWZ49pC2a8Y/Z69ML8dJqOju7ljv3
CLdkJDEh3tn1CyEErfWJ83ge5m9T8DPPxO3ctlzTh9gnrgjRqOMRtoQoqmfQNOMSJ3o1aX0eEI94
q3mc6AgX0++XyHqaeYIfFSJ9pVmY8Rxr1OA2ThuH75pm8eNxL8eGb4jVubw8IKBPKB6bYpVTutbX
6uhyNKvid9M49u05Fz1Jc8OgLBSKqgKwrBNekuRJwEnwKUmRVACPwUy2ofKP0tMtjJwzmCX+cGX4
LNtWIBCNKaQIo8SyfekAXbhPGmTR0QVXTEnnbdB2yN7xT21jO4u4uaAqOWxtja0PZCF27s5te1eW
RP977446Q1ipbORP49s6IOP6tZf5y3aO8Ujf5gWXwJEDWIEzkpQ4imlS0ybHSuJCoAKZdkStOPbs
Ekj6He9ogrP5p7Y/oNLGpXmgFHk8lyhTJEhc1HUqBP/sxeyiQk4eEUqUvTv7GxEgW9lkUU852yo2
dGCO4lHYnRE3SyhW16LxDugQ8E39WJXlPnaGzcj+/ooMJh369DoPjIOTwTLFN7uqtCA45OmRSQq1
mDq3nZhnPgku2xzdcaTtVob287wQLJb3nN/dDw5UhjJiIzptjJ2CpHVYSmui3WH0Lz/dlIIyCXaC
Ud0A+qHFLghN3oiKXmShw7T6ATfGa/x2R5neo2fuRHv9mWASxbU2dxEWViKJP+Fc2puykRp0XygE
/0tvqCaLRBAX4bnmsmSX6JGcvd1NE2+JGMFOfBnkTxWEuyIyrCq1YOwgaAvsIHXVnABhVhLwmZQc
wLH4JmOKGjA5BgKoJC/I7P/M3tnzyC3hAArTtM+Q/U3dFvW8j0psT5LSE/XjAH/1FuvEehntm5pB
pR+3SmDpW8H5qIrRgH3Y6w4sCTYT6jJA5Ve0AuT3yIQ3TM/R4eEQPBwbkRodKcI1EZnOgQa4PXz0
XGH2Vg32X6Tac3qOh4t9ijy52Xtg2AsGx3xKQuPmDf6bUmcPKxP5AgRVeZxQ627Tho2Gy+EJzlmt
bknMHZxezj99SR0094cGlMVsKISleMK88f4F9IWON8CCox3dkh0sJG3yfS/UANzptNjO8Y691uaa
Oj5/rY9HFHqL/gEwz3DWzVtzAa36VQkWglsb9cC3GT1wz870f6LiLlDLdkq8q5jP1Ye7xDpHNVvx
0DkMOJHLdE6Nl8pbG7X03V84RYA4cml/dY/JZK9eZ3NtdMIchBGNfpXFIR+7mvaLY+q0qpsYBj2g
TVzEgM0DfaTg29SqoU9pqnfr9qTCJKwdUgB+qR6o9rR0cC+z2NHDOK1uriWQ2htm3acT3SeEjjg7
a00tpajfok8Hyoy4Cm4CWagNwQoAiUUZ4363mJjaFCHvnVR7Nb5cPfqhts9oG1jNSC0hLnhhbtfD
nuRzdKgmyAWoUvpkv8cGNlMbfwEU+WTOpJOuut8IyIchQflgPZL8x2neLwhzFQ+33+M/S/Zh3sKH
+/qAsmMmWbzSj5SYWMZOPt9I01wNBjbaTsPA1HmC85x/5OO9MxUyKXTcRwCrenFioQnkzT/e7TM4
xVQpK+DnVTyVtp9X4gZ3qhbF5AltVsNxfwiiCZKT79U7bGgFewsHj58mFFZMag4Pe69bT5jfu6ww
vkzyP7tnwf4URaBufQmnvbSVjBskzb0k3aMSvvnV8F5gkeFd9kYtcc6ORdauttCtJ9wZgHFC0XpG
Uk6m6IbZPziuJ/O0hfocHceDlIe/JG/NcuUHFkWnJfv1TLWYGqcCZySq6s3R4Lp305ryRVARiGAJ
oE7xE+pO7HIJPfcRctN9U6LdSxaTb+38iR4SXWgNOaF0bIzztobA5Ap+HRHFV4wge/CPokPDG1qG
RzCSN8uRApssRk1/TSdB9hIbh9iGKqwF4xGiSGPErkYI+itmYdbOSrZVlyUkbhdolDjXEopyMHL8
eKuYqxihTNda4qcBOd1Ju2z13S7Nzc2feHxb8xYKoVLSdEsql9KXEY1t0SS/xXZuYi7aSBaoi+eY
Hf9C3t77M0fn4/lQmNwu3EayJdueAQh4DS2Xdj2249R02eUvWMqVEJQyMjsuFbTa4itYEcXbWBbX
X23h+b0KjpqA5HsuLLZ3VsqIoBY44vfkK+8CXJhPPqE1DjuTeJTqML7G8Kb6vaf+bugbOTak+CKG
WABx+DuxTm16tGCvANnukNLZUgXhm3dcDmUcVsGDLkakEv2VM8sBQ++hjCZHel7mNM/gXY5a3akt
9BBVC97SxMMm6QyZK8YRn8hj7y22oraeCjx5QuSwuy8iKeCNtN6SP3U3gHl0uwIFecERRoSkUHSt
ihUUTH7/6yPVaNElzqvocpqhXcbmIb+YPpR7ZHtecU3zKmkkmVE+bwHwnA6t7haMzj3zOqCXnH3c
roHLI+Nb6aTw9EJixqtvL4wFt2BXeMYTYH0rQLnmFhsIXzZBNqknVSk+el3+RUn03Y/oPpPOFoEV
qxg8NTQLNy98eguCdOOZ6hHX6bqKZs3q+DUFarXKOqllDJhTpaeKacOtLjNkeMQue4hMkeAyaRRF
7bKt6ejPc0MmVA9y7/N9cq+IqqGXqjXozXPa4zYr0KGpHgmAQZmqUkF/2glZGKiubolPv9apZqrM
RP/7Zwm074AhwvQVUZ861VsdquQ+QBrBHMubqKPmVCTE5jHpYOlE8Qp1y3AU1txuqkSbB3THIYEc
VsZiMSDuc02iB73Lu5oU3kyS+z36+FZEgRcssDZTPu8VQtkDwkTlgpNNEBPykO/BHnuLD1/3BlQW
X5+NjcErte9kDPOD9ABQP+A4cP2U+xHtPoPZWEGpyQm2nF1l9iYyN58GQnVyClphx03h1qzt4d+0
bjz6AkY3Q+kgRGlLL5+MU0EJmIp61CJItIBT4pkn9EGIkDnnjuHQxnyIgzsl3sTq4U8rlIuogi53
k1INkooYiRDSuvqx1OqvfPEAJ/gJBlGOzc/u7YJQovPWva0v6hthxXJYf9dyFoJ0+nD99Am4wY2D
MSfANcaaN37ALMr07KWHPaHWKDvvsYPAyyHxV6816STilikSA9cbr8nw3x6LCdMuPIbrBS2An6Jb
4xSZj0/iThKQI/iQY6ylZ63ujZvqVBrh6GTr0QGwlhFjaaQOfWLE55uDNczNiA5y6xBh8FAJDipS
HQk0SSYwHZ/yXS36XHxgkPnpVZtLFlaG7oUpQGDUG2CnY3fFKW6r1iQEgPnC08mFzDfbUFkCYORW
siNlDsJt3kWLRG+rdjHE6aONpbj17ceG/N4+Um6m3fXed0zm2Euni6yTY/M0NvzUW6aSR6ZrAPtE
mDv+AnbEEwd7APWeb2a2xenXq0/awFuoWwr//KJk32YD2MSZrQQwSuW7PSrJ7G4NzjNlVhjeXx1k
0w/vAvVva1PX1vBVcyS91pcKNFV1NS5C32Je/lCtZGbq05CTMn9TuME0qEXjmMKSxy2ju9XgJyd/
lbAYyjedh0YuDyNsQd5cCJaxwBGtMjQztTabB1zAjX7tvxIJm87VvMTIjIZKaCKNZumEMJDIvuXg
tRFllMYAdzWuowciYayA8QdMI2boCz7hr9cuNYmp/BkqxQKtOH9e2kH/Tm+VbQpFBZaXxM97r/Op
xwwbX9vfVrc7TZo0BoNPOulNB0k+KEJohtHTWWlW72Hkem0tAUYcF+8x/Y2f1FSmV4fZUADnlv2c
X3cTENmc2ZkGDmWpXUC/toyFtQPl46mnHWkTnCOMEOaTQH43TdieQMZET/XuevTofzGqZ10d9Mwu
pmcKoDFYHaqtAA1knIHOHmFO3jb0jk5D5oqMxhS5gjHFUw6mUaMbzKuabKSK8GMoSv5sQItDzL8P
hirD4LJzGX69DcCB5DI6sL27RxJdn3t0c46eiw77RrOiwNvgH7z+GgtZJLVyomBGEP/CnbuIPjwU
UF5m4xA4bjArV5pOQ4bMJQslfdQHOnlRW8PuDhVc34/lRQZlElpDkel8bdlauz8ErEw7tQ44vWjB
Tb0ZrqBRzLubzUfr+yt/28N7URVJqEJKfAh4e9OR2PHLbaE+YvWtnlrpLyBSAbzxLCoiiD36vKVk
F+8ipZRKZWWFg27YlRg0MKy6myXrA3N56vjWlZfXXMjpMrBKka4X7RHSol2W5u13pkqTdMzy4MRF
OEx9nIaeB3ikxyW/ODyxqzfp3oqL85DTl/lGuVNbIa+Qyr2OSWo4jBWnQyutZM9+t5tGwTgOL6jP
EqVN8jIXaOjnxMurK1x4fruZCsPj4pNIMHgyhtvwYkdwMV3uejjDJyd9GJQY5WINhfNYbepStuBG
XUwuDKsxyQsRpVsDu2dqCrQBIp4uEUDoucq1lyGxbuImL0TzmCFDHXkj6SMh3llFDlf2ABHuxQlk
8eCyK7k3wME9MRLMOTL5tZCVIfyeKYlQTg7J80F8G1KGQ0u+98i4ZsAcpUraVMcUXYYSBuYFwnjz
j0y1NRZRzt0XGrUsPT9Ltu7C9R0Pem+iHDQwyzlTUlytLW6P8g2MFBTKgWbzGgDOi/GOusNLjIbi
8LbyE6qIY5/hHXz7nv0qNvNdv7Y1BrUsRM+o3231I4cXEtFah7fpqq2izrR9DNEQAopltV1njVod
GBnhScT2yvXo/KS9n0wgO/ImGRkX+4vyepjyIjfoUmwkM1g6uM2Ow9TX4HPy6wBa93HI0rOOk6DJ
sp0AxTBu6fZyjxWBw5dkrlzNgDHkbLmfbwLOKrxbIRESbGYKjLkGPMN0jH7ufNEBulJQCpupp0gV
EoYKyR/FPSM6SpXd+OJ1PLYXFUbVhuxJTRixkG28uiAp+OnJywK/CCiq9lIJXKhu8U2qeaGSuBLS
HrJ0vcQm3QwlmpIJCc3jnpSaAQG4rcmLaRLdEwCaLx0YaqXkJXyLBPKPW1ECucgnKkyIgEnVBNT8
Smek494MOINyHnxtOy6cPPgQJCbbemyg7A0f/7SLsoEpmfjFnlpFu0IZPN9Xf4eYWCePp01alIZE
r4ZcBK0J59E7ALHT55mxsFlOwtPCcfrV5iT8+PEqQqrjQxoXYWv2T0JtSlLK/BNWl3P4tsOZVZs6
QXG66A1nEdJ4hX0VH5PiVgnaQANErrwfcy3XU5G9MPqxUD2KiZbFEeZxV+j5yt0XgPU9v69nS3iO
SUut4mTKpQv7sOqKWzCaL59eU92dSYWw/g5ChJPh6mJ1Gx7LErdVtfJ/hWKmeXjPCzUg8TEvgvY1
HesPvfHJi56JKQntsqfvHcORYVp9C7qAo6/YBd9fE6cjjalO+VVl8U7/z0VuIEum6b+00GL+gKws
xAv5FjkY5n024AHqIOU/B1cS+e9agYqsonYGWAmflPuOx/MIdHakWh7uEPH6SOWM06fif4Hhde8j
7B863dKMBQN8EqLtTTokPdUo4YsRElmS+JvGmdSfQNjxcIf1AxBdp1vH2ORhp6kyJRa/Cf2E2KAC
YtCEo+I6SgBzckqiWLIytgocXevkPr803EZi8nzNJdfzJ1uce0hw4Xg5tneb4lPM+nesOd7Z/m/E
Gysyx2ChYdfFIzEb/0GXzBlSEkCpwptv40b7Npx9oEnrt22CQ04uoRMX4l3QzI9RqODPod0qjgre
xAKXZKPRN2rAQrRN9Ortqq4ZtS7TvUKpGayU8OQjX/91O/zFRkRLc1mhFWdrYhiPWEQn3j06SzKB
sjKWT9mUiN5Y4t7o60LHinmEzk+Se+G7W+PPsszDUTweZiEecnYv9KdnLt83BO/xpVVQwzmzbl0K
ZI8z7hsO8txXlCxP/yEoBrZjE4o0O3zWagaVALgcxqv4Cjx4MNrGnNxPu+yoIasQQjZ3TXfE6DoB
NkMP4EeDSnt1/z5h4Dxmxe7h3vunwRtsVPVmDf/UGFgr77okW2SlZs16DLxXUjn9moD2oF8Wzs+t
yUAUsNHurCW8j/yXBX5XgpnTxrxejB2vbnFl696EvGmvrSRnIE50EVWQeyzEaoiGxOVDoap5Dy/r
ssSmryEjmPHesGwas2v5+QGI5AureUp8YBOSy+99DSqecRdbDfMn3zCh3o1xQsHqXXD2eAnSdyCP
QQVqLrMLFTR/PXIpjuUzH8xp/z4ioaiYxLQyPHjBA++Qg+i7yxD6SsB+jA5crpg1OqqaXdozn2rq
s4mM8WsMdX7716Li6U0g1W4cWv0Ddnbc605hePsVIlmzBNk1kW9LhbiqAjKZ+dAAiOvgywxnY5IO
eBUUQ3dr1VqGYpK4ZI0fR9JOEsiZlyTNxg8TdaiHfufs5TQJ2ai322yyya6gi/CrUpiMf/Oc4sgg
qn+afIlCOJjBaMRexokLYyTGkV6l+JuFo9owk/4lIkxC+J3ercIaUCHtNamlI2AyyzXCnRXkr0Yd
H9LFvXbXtR44YHu4XZFii0uWteDMH1iZ22xa3coTDCd6pOexOXnWGWSNCr4Htdny8GJY03cWmxny
1zazY1QgPh7t+rrK0DzFdc7RMiM6tyl95+mQpemYjKl1CRFBAEXi7moG7jRF0nnSsZHKU9f/o/OJ
klYqL33E+FngzW1tTjU6bta5ogxW4wOKbwyMZN15LBqh0qoZG0OVNYKegKGAekcWH+3EqWcPGcUl
S6pW7H/zKf91gIXLF85a+loD1WnOPPvZhHrjCPoC15y8msjCvT/ykbMQ3rHbxymZ/aTC21Hsq/LI
wsAK46LD7NuGf7CMSZQ+qNuU8vIsnOWB8JZfmmQm5r1Ckg4AiPajauktLSfa2xJtLPBr45IQHmRr
3SJMRHqTGq3tGUOWVHuzCs2vfJhAAPsnF4umTIT0X8Thyln6SI6WwnAjguKp4yI7xjIz0BbMoruM
L+pedNgpGU0fI9oICZLWT3yyRxBY5qWahy8SCIKBbiVIa09llBkDoIsQQeWtFyf0hxpDYnAx08Ei
SAiTnjfjgQW0Z023LMYZHJFQGgjQ6d4nZgu+/n2zI9iOlYq9cnMSrijvy/njwmQKVqgczEjSkWNF
J4azfCv03mPVYUz7+7sA1o7d1cZFFvU8dwOfJunOQBhrETj96JVX51vd/2H1ue3G5a9/La7aiYej
k1FC2mKlIp97VEoouHco414QdwtMHu7JSR0wNnS9ov6n/HfoLF3djdi7c0RqmSsULyIcWJDcWGDK
x8pCvqnEjOZP4eMToPTGKtBZ0Lh2QTGA7gWbcfqFrAuZdI2J8Tmskf57Pz57fW7zYlTvfxyTZNM1
YLnV/GBv2y0OriscqiQmYUPtd4KM25cRf3IF2+xrriOoc7M2s5h3/bZSUllhhR60pzqpHDLsCRVr
MkxNYg5hr5AoYSJkDPM4TE/mgFsTZfKViBDI+1JLb8/r842V4vFqYtafsRwp0fpdlSzTAU2TA73e
h44YVvNnqKWw3XmpGNMrcEJ/cPmXVfoHP9JWNeQAlrfg/CV8cHgJmB6d/QnJjYgIrzlhSFCjaxk2
xEuKElCuDDSQLRGZ6/qny4oxCJUu5A/eUiDMj8JcLdeeqquyvPU4G8ZQzW1WEbJehsZWulQrZvJ+
pwY+TY/LRzyMQRvmMWT4p5DXLLjLw6tJ2ZBHMw3z91T+CtCcKH3hI5KUE5iV7NGdp3TQFtYut4/X
P0le+7pmAI7NbC0+yuWCBdfxoqY5rMt54XxEduQMLlN8w0P8T5MJiyGPbGx+cslxUmGF50UQ7MWt
GNTaDLNqpCJzzWVzUgJnv4cdYeGqvey58T4z6OwU40IvGHwpzi0Iq5XVm2Hxr2NgrpkdcShTrchQ
rjM3NjN7VqRz4LMCPBEW1IgRMC+5JTnHkyp06XOuDPndcjblqYPkgcdxUpEDjp4IYmdXdz4G7uOO
7BxXIhwzxrfY4QFzEEUYnNyWY3GhEViBHQPTtLtpO7lCJ5EUhG5sExYCN9s27VK//gT2L8xa5yJ8
OroqjQbo3fV+rg3tg8vYsbC3YWtKFuKFQTIwsxXmuMh3SzHWziPSFt79jDDM8POdIPXk4DaSAfTk
H+FCLZexHs3VZwgaYTZi2jNvAP3qy5GY+3GCAIYsXeF8shuSS6Mg7EPI+e2YyKXLX0qlloQ36rUu
PHDkc9FslMFm/4mdU4px7pOppOoG1yuxSuFNJD38zUqbKkkc6oJNqcf5GJpaISYUMqcX6z4Np7Wb
kCSjaRimMXEwCtEQ/AIA2l3yt7XvjHR+ura3hQpjKaUNtIkpsKOstGC+O3wFrdBRHWJZKxD9KgNT
s6uo+MpRTsDY1ehkByq+7rtl/iB7qc+xFSq8lpF8oi7WP/BV04/6nqoad7FyrG/1/RSIoQr7pOA7
qkbGY30PQlCu0StrTGYH5f0WRrTfrYdMNYFhagNEJ0ciOmIlC+N7kOshcV4z7UKHkv4cEFdq1Fw9
toXy9fzJquCrmXgQtmKuVyQyDEFK6eV26oFvl/a76lcdVoC4aSi/SFPADa5fe9P13OxDNHAxh36H
Op+M+xtEmagRyHpKbSRTt5E11alG6mr2RfnXymKbW5gDYjp1zz8rWfYZCxEcGQvWtYTTscEOjgBi
W2JcHfLnIhVXwEXZF8ra/FJBXYxfeL2S+4Hr51IbbFJw+N00z/gQvo1QKyLyguhaqIvEOU+dZSew
omPn9Fywu9VHVaE5hvtyGwvA404tBRi8gqo3VOAY2ZeOSbslDLCJREYoZM4SGj/R/Vbh7WNPMAwD
Y+JEPZEb9MijOGXE1VKNqR01OSc3pCh95XQc/hCwkwiDA59da9lIPFjwZRyvceZFTXncn6YAmiVJ
0AZNOD5RzJAtN5MMjrmch4cCGiRoIqR6AKFmrQO9cvWDX1CXZK971x7n51ztMR01TcyflReJaVuz
zAJx6M8t99RRKDr//t6qF+Oz2amScy2Y/kivH87S7O43nohc0BGvFAAIpfr03TMDpg6omRrF9Xds
ocyg8pM2SgmH8JNr563ar+AgYU/zunS+V6rSDfRGozGJa0aglRIPrgZGe9H+QxNK4DMUEPjXg0v5
fE+woBPyC2s7ysH1rN98hFN9fVZ1kCttnRxhTaUXgLEWJ58tHxgS9yreaxFKKJop4VhH8AoXhCcL
upsMRC9TYHxL82Xa+bGjSCwkU+8tqg1jb6DTEBD2QXb1SrIO8l/pdq8G8YpSJMGvbVduhusp2iUp
KeliepRA0g/1D4bimn7b8XEtMXA5jUpnaKaBdvjmO0iTXgDF/UF4NbgvnpxNgefacJGjVC9/QMWq
tEQIohYMiF1uzntvkV77cPITVrNtAjUPFALnH0pJfweCaURjbTX13reV8FZJoGoSpvf/Qpm/TxBx
cxGGvtOi5pRXRcQtwxj9/EEDYpTT/XJccKEdSD7JEkCqrNg8izsO9atpYfX9zDiHXt6FiaeJrYJe
hRSXLFTMPeQLv1C/V3qXGDqvqEasZom40ocqiFg31Xwn9PqFTpb+gVX5UY+PennbESlaVh3/Z4UB
JDWBVu6rZSIETktaWvgB595ybr2cwQWPGXg9Dr2LJRNdCZnauzH6VwgheTP1TBAa00lYnid6vvZi
I5ZZg4mutqg315nQkKsjkJf9UovCcuF7X8W7318GaIQW/6sTHzSKywpYEIw2WXss0IOayO7IPwCV
LTtNQWwCu+VN3q7RLAnReuWxwONAKGWpYsZ+2gkxFiWsWeVxPX0fku+Qt8o2cjx3qdG4BObmqieZ
Ntv3TwWDZMvF3ySDhFpVA9ZyrvqafWiYZtkH53FSLFq2IpGfjNCGoF/QYZoGxyx5mIIGQ9L9dk/d
FdMubySMsqM0xDOL8D6JdpFg4Gn+UYOBZ2G0So0J4C676EGgq2+Ck58dBGZQa8DefqxNw5qOwzIV
X8Q0x0JikWA3o09lj41gxzW9VktN6U9tN5g9sYFNZz8vyFvMH8mqSYbMl5yPulubVa4rhlGCMXKB
NiYL30aVLul+dS5HFJRqQmGrJVyvVmppdELW0S8GCgtYYQpPjExiAuGNt4nWRsquU6zv2ukBMTMe
SiJbvhB7TUKTk3+bqdcB17hccSYdssgl45OhtrErRMsWeMuNKlMvZ1KicYGUBNtAXPbxe8WTozPW
YKP+QVNjRGVAu8xMJ9xDGYBkQfjAWZADAdKdE5TCaZII0bt4OEcCw8tFS9dGK14HxDZ9eNMbRHXL
p+Xv3/9k7NsNHxlWnKsb891Tj6dgqH6eUrdzk5D3TJUd1N/UJ+pD5bcu9yhxcvZ669qEr3GXdqDS
Ui/RqJD4ZQEyYcor5IzA94FZjqL/qPX2DxroADUdrbR8nVFEK0oe/ZSn/+jRaaKaNT1S5XMJaia3
FBOtXhwR/bydwGekRMYs3BKqa7ugdraOSI35TOkzEyvnebEW0PLGui73XP2oxdJxguKpgTRJzB4A
PiLusjBCMKJBMQxb/f7gDbDZxYA8AfxYeRsIZv4Tun71IW2Pm79y8pIRrJp63mT6seLP+fhkJZCh
+jqSlE9+PrbGtwWG7RduAxvCH4hlA/BBybCgS4k2x0PoURxAmEVWDk+Jc79iX3YqPCjyAvDn7hpy
35O+/tcXh36xcOTor9D3JsRTwJwmCLCpemUOczm/cZ4IKfv6eng3rhUA1rax6U6TLiNZckZeoGuJ
D/F2fAaZVrKmpnbbiv2zN8mnoKVVBuWYVChcBncu2p0M5UzYEgtGqvpEV/lHVjJBUX8ydWLvK/Hf
Gm2gdvH+0xkLFeluXH2mSJliwsyey+pTbPS4Wy1Mzq31jf7Yb/oFKzWSo4IKera/KUq6kP8n6haF
mTjs2G3xVdFo9/7xLnbAXfbR+p4Fgyy+YQersfkN79Io0akljpa23HiMq/bKAeY6rbLnY+BnnAXz
DVTgDSN90SAWlcO+JJE49Bu9isIgJUmwTPxXEPYkR6ecmcwk5Nkr02S8VP1gS05fJvoDTliPgP5h
2YTkQL1swUGLk2shARsrIP8VXQ9Kt5OiEF9XfgQD1A2AqlxREqqAl2XfbuWyC2wWGGLiBu9yp7Fm
uR8QNOEwlbxv5DfnceaLX05qvllrFmHID14bYVe43fAUS4p9gMLjQdOR3PmE4DZ+sppludxXznQc
MzXfibaSFaNpuj29XuK8n9ZpRIQ0hV5N+k9Rt5nmIsfSKro7gpGaEOmZx3gG7Yyks1UiIgSv4RCl
F0gkTqOty3F6MAwjDmSzEDZJ0DowJNPH29ex/efBZPAECtE70V6BAk64Z1w4Q6hvQ/HUcR4BNDjM
v/zavwYXRpqMp+k/oDCNOQ6bV725nTzkrfX1greQwX/Ye7u+BdhnBk9W8+pgNeQqG8a21dCQeGFy
kHnbD/GxiTZZ6wc5XOXIZf5bmuoZRedhj5b9+BcyR9EoFgljyhBe9wqIcQCJufYJpRWNh8aDAVIP
JVM2cBBQ+Wo72UOqlAtA/TbhH5jveIrTVN+6/9kXrTZEgppdIp47PfpDInqBcsR9TmW14qdc2IUh
wnG3BxR5FAAAN+rxoxitof0T7OJVsXTzB1/NRex28lFybDEJvWh/jrLdoys05sM23bMzpPjdB8IX
XvMHFYvue3bwsV5vcQHc0LD8j7B5XDAuEoZxSYp1WLQut/kVbLIe37hNqi6Cv0hFEyAuRDQ9vkIQ
1iUmVkmdBGqZCKgb/b0fQh1qbiShWurX3CV+chAEm7ZjMaDHdWU1AINbbNclCIgwtGPwS29njYnw
AI0h/LO8wpHZHt2uxj6NTs4KxscoW6Qi4LxYfnnVM8dNryyVSPGs3CR7h64EHUtybRCt8Gu2st9y
IrdVjH9NYplWo7TvwwTjWqckj6Z/0P2TEasF9K7BwZbOdYjZEUukJzfGoY89+DsfOxEqenbW0IMf
GlZYszg7CL3SZGnIg/Mx0qUIG+dFXJA8uLA9DpznY8BBwofFC63e+zzEKf6dfnKHh/t4EgBi5x0m
uh6bQaVrQ77cuqSsiHo813WL7ReyO6UCdFA1///lMpKZksZQK1A0nadtoG0q3sn9FCX2Ifm3jO4e
hSmh+j+oujjZ22F/kMyEtfS8x3C9WeEovV4YClGzVjE3BCxyl8YO3ZqRROeelDfJaw6scsH+rpm2
mfmlGA5dmk18NdC6PI5gX4f2oRPTwXb2IzsiPcH032XWOXO3fanrZogmSLfj51r9oQ24qCR3z7HJ
eXNIXuwOaeDO4Zl5U5TT9kLe++Vk47nqaKlXW7xvPpCRD3SnDGD3lJZq83v0PXBd9R3QPupYmCv+
2u3aNppKwL/0kpwFNy5NqST5iQ0pRzjuUaK1SCYfl4M6zhrKVjGtD9In9FGGrsDDQEVcOhaHmcIy
3wiDoI6tfuxBNxEvYP6pJJITTMXOGu6L2KG51Vy+9iVPJ/kVmIe94wg53EFVJyFOwvCwUg6PACKK
w3CcXknH2ho+lSgd7ouwM1sUWKe87Y2YXt/FXU0fuBoFV9qgyv2LbTRyrSqDpxQNlJZcpCPTAejN
boL5mzZimkMssJoCU6Nj/6kP4MrF55K1Lu58hRGM9NbtMx/uOBUaja+mcUS2YTkTnmxuGGibfVcq
+lmpLxtZdtEPEYG0XiMzPP9Y72jp8N93gwyPGzeVFKkQ4ErcXG4awSsDg8Zef2R1OlPMYg8fgJe/
7qz0uGP9YsbuVb9w2R1LNyUNzbVqYAhB1T8W2PhqmVWaP0BOMbvFTX8p6cAzjlj2fsh6hoekgRdz
489Lq0b5+8nl8fQ23XcYl3/d37AO6xofpwMTvalPa5E68PkR2JCjcNL+yj0rKE8qiRBN6vvPyCiz
aZub2W2B1reSao1+7JtlpaH+/lnZciJJ08Qq5I70wDmVgg7XUyCluj3ng9Eb9yVbWF2qGhd/Uj85
1xufZ6yQNt/43SBPKyYhXpxbQM+Y8858VGmmfVmZqKO1yx1/hRF8Sfrr/TUb3h5bUg+sJZPz/Y5c
EjbHyNF64Am09XgdQH5u/L3l58AsutZSaxwHKwnlR3uHjj/shZj+kQmGW68xFwOTvIetJINZkr9t
czkINxKJ7r2P5okBJ4smSRcOkxAoZYuX5W3+AnF5Siayeb1unz+EG8fYGXVeuv4pCIdLuRhLRRHb
W/Z95sNCXAXFhX6dzEIA2wsD0xInrHXXqlmuN0NYvrlkSWFq2b1wZQOIx3HZ8WagfT5IiXjKDhdm
331lys/+sIEJ3GEFXSNwnURxp3I81F9cZ0nNhqWVT6cdF80Lof8bhO/2PyJNNhssY5+UJQtDd6hE
jufU/x1O4lO1mhXrXPApkbiGSQjJ6OrlH2+HTWa/vWg4aUtTO4jiOY+XzMyZaalO2pJpG6TUEtkZ
+S2VSInF7vZhrmk2PwtlIkdfMAkXsHHBLQQfEfUN51U8tyqidub7dc+m3zKs7I+x63u82zSxRS5/
Ani/vDJz6wwd2MGAGtasfSERWMvPqZtGGgUEIA/tdOGOnf6DIKIvKMGiBDG8QnBsIKFkIcxB/7YB
sXrXgzkrpa4L6yP9VP4LLgZ+erdED97Y3yBAp6MCHAR21inRo+GxfJtA1uwGpcx1Rmsi5DOE9LBv
GJhQEwNcuU5ZM+6b46MvyhGKQaScqtP8s5JWa0euJuGFwXl2KyxM4y4ZvNG8FkMBpQrmTBpS6nXn
TKm6CY/prlDkJBWaV/ZZq28jKtW0N8lW0l/bENf6N8p7rN3xk8jLbIbM/YhCOocxjXm+hOQOU389
EqhzUYH2prNkR7Ckrf0GP3vukywd7/VlZ0a38IdFHvcjdTRsqbhDovcHwe8t55xBGEIQ+2frk6Ja
4d59m9uyj8p7HkgMb5bPPpov3uoWiNMwsoaopjAO+xqDHy2QTJj91A44Ee7c762aBgwr+ktBCZmt
6smti4QhdWE3DGDdT+ekdVf2t2Rt5MIl/sfTyuWV7As7126PXkotnnpSr8/hto0P74/ztHMiHl2p
feSK+4JmzfBjRQ8LZp2sYcQimuJHMxabmzesbe7Ro6EQgePFciovTIY2MNCoDYyBuTJGfOt/JZ81
Ysqj2qLYpf/jQawYpmcLRqJEF6IqreBVd67ICV2P9I4slWYOu/eION+x6SWJFbfDQUpPhuCmhPBs
+uiDf9ENWiSuujBFUiVsPKWW5REqJL9JWmoQ77rXhPkH8Oa12O4gurPwkwugarWsnJTNLYlgM8Ey
FLaoxK5knFZ4uDOdVRv34U2OEImOyMaXkD286KhpwG5IUrNTyRdesybT4WrR/nmZtn4CaH9MYGpv
vByOA26+g3SsKZNV3eEEx+0mk78V0kOSlkHeywTSFLyIzCH3zUWQc+bpJz8hAgJmdYeF5elzIhkR
IJfEHOGJibrVX5wd32NSnE5PKxPY6UBcgHEOOi44ITOqtsK31sNY7llNXWtKyB1iq1Fn+pHO2IwZ
wOaAFhd3JUBhfpniwny/rKPBr2tCfeEv1zikGK3edx9aswRxTHxnypWtb9D7rS8qm8rsmsRjSqT7
9I6vR6YsRWXP9+frNI6qdTSGSzLaTJzB1RUv++TgSlPJ7zAzJc+AqVNhdOV432Ys8aErGU1oXHRJ
RgmOSsjyw8Iubg5TDnPPcHLYVtbM7qWv54C4cXoab8RVSbxJ+KDvHRWEj6hOIKWAQZU3DlEIzIEm
UyXmGRHHz9L3PxMViB2rBmICOkX93vFQgA+g79rgebv8a2PGvgFKVr2l1VrWPL7Fb5/Glh/eXkGX
FLIhf+GuQYNVXYWNlOENIkhDZDO8fsFeyujSqFREfgRp7VD3REL/HSGwVxRORRdfZhtK8SiBsVbS
hX8DY0v++6y+XQ2hAXHXeb8HBrl1kDkYpef5lvT1lLqv1yoUv1pxVjz6wIjGgCZnT/pKLJJKFprJ
edsetJbVm1OhrmepgEnuIP7LVKYAUHlkrEHWP5GkYBgGWacJLNwv5GwPFbtODvtoRtAi35dppIVu
zrnMQNi/zylLuQZudn6Jgp96uHeklzXf+VsozC+na9LQZ4bDci3yarB6G0mY2UWtTAM0Tz2DiDEf
cUHUnQAm22HgYV7DGblMBSajAdinIVTBlmJBkGEJFSFeUAJVgrcYc6Fu0hauuxvHmZ7Pg4vbNLG+
gnJ3UxnRoLHXfkh8Ll8tE8TVLq0UwqbkEEHuTX6WclyRdb3nKYQj6U4AFw+YLffNBDeXtOrL809X
eSLODQBkWK5odPtY/O9boUdDdnsEKuGPXTrbBgyj0azIdkEgaVfW48oi77Ag6cRUI4AIBbY8iCi4
MCxbeFf53vlWnczkgcrwQ9q0SwgwBkzEVhSDx1DBGjBoq6RFrN+3uUc+/68nSDDSN5zWMcDmQ8Q9
1NgQ0OYud4ZhRHkfRnVr7yIB4tIjyOh9tzum2z5qeMzTGaSBGx5VpUPzAX3A+ZblzDOelwfGbcoK
mn9Fx/5uz5xw+xM/eegoX6ROTgO6tecMn49xQpJJPnR8ZuEIfu3KmZRmUho1EiEudZg/4KN7HDnV
aqkiU2kKggft2cbyE0+ll93WBhEXo9Dn2TLmgAEn6wmyX65sZXGUXdlMjjpnQtFevoazJXkygwvZ
OQxwlPsI47BRvGuxLi+7UGI1xEvbEoZqIHA+/c4klHsVGVLRvd5zCq+BD3VzaXqaVzrZNTPb+w2K
YDQ6yQNE1gTkA/EUe0p7cmdHRBi2SJ5GVhzkxdODPrvajr9A0g60VdLKXQ5e8YTloJUgBL3MwQlp
6YhxnKk9bkmtQuCxBcKB3Hc5c9wMuc/BPi8gDJDBUBcCjCTGiW3wtLigOK8Db7edHYJVSOc62sb+
fQAZARgTHHHBVfyCVKNfDr7TWrV2Z+zFliCEKycLDHQYjETnI2yeszLCHfqap7eAJVzgpNxyeWo9
VwAVP/QSekeD2yGV4fVgMX8k30IuQ3S1q50B11dXsgtYyVVMzTWGV5bs8hg9dDQ84TwKArCprWwC
65Ms8ZxgnAkDvS5LI7wRDSrSgYxLfMGGpmQJAIDWqS38spjPZI79CQseSWPSgGQ6rTapJAaV6FxN
96gEAiC6NSOpqm9dzQc7oq4u/SD4WR4UUZD0jvyzCVMAdd6EWV13aAygPw5iQN/R9djolOLgewUG
hNzaHbRc30YzmNsH/jg3qqwB3dZDIAUBPhs0fI4fWRYyQ+LA39mVCN21kA5fyxPvwXdyZoXq+2sX
gW8liqK510iAI8TC7Efcdgc+iBwbtjUlTA572OkXz1Wj4C1CYaTwMTxo5MLoulG62PJOfUdtwcvo
ooBcMA+SYHcftHN7tZGvq33Jeva+LQeNC1e08saaqnsUK746VD0kL1RUcwGxvQ/pCA4KI0aqX6zp
J0TysziM/mFZ/TaUpGrXHYxl/SFPVFnn9tZfhwqn25q6dG3nCKh7SFVY6d3beUX/2TmjCEXL/nCN
3XhrvJKretHzwvt85A7HsVxJoOrmMS+iDTIHsnL7ElEoY/v5ciN4LBCEEcC1Ufx0Q7hFid9CEO0r
/ySwKal540qxbqlqprXhw8+Es4pX887HasTl4pvwLamm8mJOC/i8wMsdu6I7xlzCVVHQNjvJ2NYa
Y5L1YwxN0Opz1eHToYTxUX3KJVRw/Xd0B2aGZNjStw7eNwnuszHaFUN1+D0eKHOYScEsnpD3vOUn
tVhwelNYFf3k8wdBSmdRyocUhoSZf50lQbbavMZrYCJpSbCi/SGRyR3sQRLXoBFAuNP/ZzaF0Ys7
1kworVaUkcOXorGF/2WP9CJr9TtzvA3XorphpK3iSO9Y3RkrU1CXHnx866Yh47PLGzk4JiOONyzY
4TYQnpcLql01hwpFmD+6mOoSYIUoJ0K/Lte93GBCJKuql0DGt2QueeHu5VOn4yB1Q4gIybGndAnE
7dmytHgNbLj+9gQdhK4MnqUPoseMlzG8E/kzQNpA257WlJ9yHmKavl/R8M8af7YdWYO8O/TE4Qwa
AnoahBbbP8SOHmDNPx0fObWlQ3Oqpq53G4XuRlUY9KZfZkPBgBbC9UykeYXUx3A+NIKzETu/s60N
Z5FX62ZJvp0q4yoLhOijGrikCQx5QHnb5k6ilTk38WvN+9AnfsQrIR3fqZO4zFbCLa+O8eR/fYXo
yTNt8vJZGbcZeqacd369bw2B4VR/OejYRuUnSZLNoKzHjAQ5NT/mmvUAH7dyGgXRcx/lSIib9rxG
kiz8KnwCtoUX9njIeln5h+m8hkRchXpi6VawlH6dq8x3KpOV7fwv8xohKOGGdqhTeoCm6fSU8lYk
L0IdE3RmTZt/cOADLPE4ZtLJPDoH0m3hFOdUwAub740AwMeq68JJtdrTA8y3LHAmgpScjmDFYq9A
bH8y2DzN3kEmnxg40bhBdO8u5ucXbks0W9+6ybin15uq50syPSUbewQGYb2tzz5h1fv4PsLXkWM/
5oXcbUhc6w9mRxdWOTe0XYAwHFcH3dzo9lPmOpeRgLhTDMq8zV5sSuZF3IMpJNrorWcQ4xbVC/Pw
V7uxGwY9MxjKf6Qj7Mpas7MwiIrqx8Rt8xPnyEnyqybFzLAOf6GUBcegPcvRedNUzN3+5SycDNG2
wbhj6RFp5QL0/8Xc3MxhmSHpDTUSosfBIKbxi+pxvhZdUB672Yv8BUc2LJl9OQxl5f2n7zJ1FR2J
wgPMSSQ/3XYES5ZR/m7NQHVk2xVznlryJKzsjFdCFwoa5PV7Pw2BxNFDzaCj4e0Fg27yErnF1dD/
mbqvR/BCzDVPr/j6wQbMTBztKZxuV+jZERiNYLt+PPnseDz+bv1MIYBVmagNcNDwVsa58n7rIctf
pbUI80koTY6EeQxihnb45J1W3MtMge9gWnBkVJM4AB3bQCAdRR0ewlCSSGDc53FHfH3pOe5PGDdG
ruuWomywXK7IauPfnA8R/ATBO8bub9MtjNq8wVdoB8Yb3wgHOiqfvHPhrcvFr7LqpOf1zUnLeQh0
38ZSPbILqaLiIeAXRd5cYFfbwoVtEJ/Bj6meDTTIsBJhbwAwPG/r0PgU1D8fiNQItv8u01vMJfU1
Q0XBiQuZc6CitzU5dYogAxZaiwxmb66eJfze1Cdo1Ei3HNDbcwRKj5ClNQpffERUI9t1+bW87Njf
fssEcpLlZUcC8FqHL+BW3UAxuFNZZypBXUaFRjHB1AwybkDhUH0HZPuiF4FRKJwEvwiXHlLdH6IN
Zf3TvMSzckm77KPpxmDe5Smma3sTCMf5NH6de1cNZ0QGjbMwMgd+hqpWPTGuU/bZG5dtuj/5bDhy
s2nwxod07CqxDA7o0RynVNFDee6M4hcwKN+k2hPv5d9gimp/zGki5EJMLXl3TGeW4Cl9HVjEYYFb
pbbEl47DWmlB1KcoZV7+wyrPatg0esXBB7DBMUUFP58DrF9hkphgsX4jjEsVaI3A5isFhTnSP03h
CZRPUMkFI/5gbG8K0EpHTiFZmzANBTW0hv+y7yqDIP/TCwjfW92+UNJhmr3H5oqUkO8cXsR1M9PZ
8JZSgyl5hM8+RelVHERnCbmaycvlPxfQoEEQcxFlaVMkabx49RuSUbecvspYcalN+ajGC6UEePTl
ylj4JyRggku9JlAIsrENgSkq6COfcVd8QPvbbLvRCnvtD4EPOxS8fv2OMdTz8pMypfwNU0IMsA0u
Hi6x0bxT91PW0LxrwVNCTsNikP8Cb1wbMEqCulGXYLqLP9u4dcGePpmu9RgcSqc408GHlWg8Mo9A
mLkCsLt9KfhLy0STWgiNEiT7cGGF05AeAO//5ls52DcjxqBP2zaQmaPkWJEuYzlPLvJclH5tNlbV
QcAvBpo7e/YI7e4Bek1FMtneFQ00YEd3qnogh3zIfNigBLyrTjFowOcEAz7KjZASmuHpCTYxq9Rb
OS4zE/NnjCw5OqRE+qipdAEBN+W9RlSnhyazuM7xn0r6+Eyot0oQDZuUXNmZ9H5rztQ0kPq78ZfT
escIF5IO1YrsNS7tFdc/oO+hWKbXrhAHK47EKSKv3AoroEBXLhFZARO3vAaZVldrNWZhzjq3TIgW
Xak2Z7JGj0GrIy/xR8x79SkMlPj6XqVVRRWjjfvv4dRCzw9DNS3rALPYwIkvz39uKx7FmS7SY0SO
MyTlkX3Sk1GWUYtS4w6+NQ41TIGjChaG5MEeQ0hWIWwsvr9ydmSBit1ItQ/YaSKDyLlKdpWsZ9ZR
KQFqeoXeb4xc10qP8RGbyxupmrfnxn7J7e+7N6Pcmd4ZBgYZr+L9LqZHhW4d4maybgBxYUCK9Su+
6sJuo+B/HCFCrtgcqF9eY+FSvh2LeNlpI/iRZjiWs4wPscOi3yJFnwgpFvReFGY51CRf44x3x0eH
4Ee9K582jDuIACgiGD9koAXV8//swXHG4l5ZU96ZGARr5dROPva2vWL50bh+0ERArc4f3pdDb5im
QtH6lxJKd32prqfAsdLis78Zs5YZaP/GHO7EhXdGVKMAeDHvOooglIVk6UoW1zXR2OyW9mC8nSLS
ca50Whxpg6NbdlbtxPVPJA15veZXiu+6NzwybrDsbtmxHmCaiqlot/pCjwFbkkdva6+Al8qBqCF/
rC0DsTX1pwyfo6RFIBvvfuWiGjwDH0AQYpllubpu5Y5Gd6x/NzFIAAguM6SWTbWardTJOyUQO5Ip
uVfPC/c7zf9eJNqddMeoIQUyh5+cegjSdQk7vb5gI6k10Zn2LWSPyy8Odp3VEKR2ZFXiUxQLt67Y
c3NyXtQDHYnF6DvmGngPEG4hLInYYw9ooe35k+xJoG9YbRwlmVYMwwp5muP8/QrNq6+txcialGY4
YbKDmz6JIPHshrJBxm6gYGdesQjbWK7wIU94/WGFVFRFt6kpMereqOnMJbrnmIx9J2ukpWgjhhgd
IFQUAnvIEvYw6LqBwRJhdjYeOT4cv4KUOI9LiWIomJJYGNyQ6z8CFtkA8Mwu+ltxBxHZVdI5sXjj
jXKXDyDf0y57AUT1xO5KwkFhAE0DjNKHjKBBckyvA3wcRAyNurVyGLvNCdTw+qPjRzyaQUP9zlSM
abLmyw3kn93hcFlWY3o9nYXX9+m9nVNqso3vqn+bKwnbttdsvQeucKRVqI49oC6/5msTcbGRsNv4
BQq9mcEZVURUWXFI+pWgKIq+dzR4T8QfZZ17WPVnEbjPKdY5u7WFFIyAy5qoZU6lSRxbCINsdgKl
moD/GHX7cL8pBQFZ7cbA3cYOgejK5pLHjVxJI4pKYyJYhzz5Djbv8Atgo17bzt7ZnUa2FVnPuEXP
ohPpuaSCgFj16SfZ3o+NcO8SkRq0poHXVNgkqWxrAIDNuP9H7KogqNyFrZHCAgXA0gEp8Vp00USY
Jv9Ipf9jQ/71QdRqCNonizjonFFc6JlpxqqTIN46gkIbPHi/4H2owBbtUo4A+fGm+B7bRiyiauVp
rhpN/1gf4KC4rbntEtfuZITtszJ+NoVS1M8LaaMIF3pQOIjDxT6+IDyIk/0MNKduy9sAF2eI+0xs
q6Q46CiUlbJ9epyMCIJVDM3sIkySslsifgBFArSaPVmNED3ckqZvkXC2PaRmR5wXDhSEl7+vsJT2
syx3//P7T5otzVdIKk8LLpn+2s5UAK/9bSgbCrk+zUk1ObY1XNYCg+992g/dlvBGhs4KJnl3Eil7
e00uhNLQehHzk511IKqeigfs70yB4my1C+04AM4uWVvsor+yY9EnKJSxjKHSoV596iIzcVhCLeo2
A69vNEVqR2AZ3IehROJE3aHM/9rCXJ4j8v8x6NB4lzJ/NBtVucm48peyWRUnpiudWMS+PfDBqVaY
YQFN+vkDBaiG3DF2HTvSeo+Bl7whm59O8DOJ7W4LnLzi/VjwW13L7bmL/K2Ju4p+SKr0KcbjkIhw
O2PCxV/Fdv3DzXowoP/MLwaxIqgrMUU4a7dB4wAXoJHY6dtGYdXVQupT6RhgvLTPV/FyMiEYvNPO
H12OQFZ1dzfvc4vJ3UpDS0pEgENETUGS7E7/HNg1Gaku6SM716VLyhP5rz1TJLizCs0oooEUyWMD
exckOjorcnDRjGqgbWVUlBHhtI1tg1ZPSmK9KmGZ8a+KgvaEEz6G0WskKv6DrVyPnMptFg47XW74
FzJeK/h1AAxLhFlyAiBx6BMbRkU+Ilas/VeUEas2QhFlxRkFf7dDzEEKGsznZdH6FtpwVTd0mXxh
qvpOla4ajjBJqhtQm6Sb5GnxT1PdPsRF70uwYkZA0sZ0mqUdo4+gP90yCsOcnUjSymr8oeIIpooE
WxRsin56cbx9DCb6OVSg+VPlbwQyZ62bIgzzFWq+RqJ2nn+gaXzS7jv3x2O/BS6uERbip0WPPQXl
SMQzpZ9wD1xXsDtTLzCrLSU4FipnT6Smv/OWfXA1yLWCqXfmF7Nt3iI4kGdLRqNtPGaL/AqpJLEs
X5mLTMs0G6hCOdDZXNT8RvnIgsZ50hvblV2foBv6Y8ZIVsYNsVj0VUOqba9FFHAoeea4/DFssqF/
FRC9vMJiz/b3WByOF6trrXGPR212rio8Abo59Rbe9EjEV9oEsi9hYYiEd8R9B0FUgjNzwjDkQulM
IsI2Mjfzc3f7fhecloaTPG/E2vZdoa9MiGT8XN862wvlK4srrNz0lwbJlr1I96KALHSaOITySIU0
5axMx2QopCX1DUrghvI6tk4ZhkKM4qZVekQm5ZaPhLAXeE6BS4Fe2VEIsqTzWol8Cq6uqDPDX9Kd
CC+65sILFi9326Vlb2J6m3gT9wC+7Xv6Ps8sPhKmbM4mZqA75x3k1AR7PCY1QHe9Wco2Bi35eQmH
Y+wBbp3lMHOJDecRVyvhbdxV0fDljVPm5vIIUbc45L0aUFfsk1wtgV2+ER7/tJ9zRCcA5y+YDllW
8mmWDy1h07kAqFUg0NF8hmVtKLMasXvg0Y9eJF8ivmWtKMd3DnBfBWb8pKo9NdjrJUKnqStAvGvA
3E9TEs1Cv+DNiV0au0ZuGJH+HLYz5p+62/i8VEXPKRAZalAId1kJEGcgSYAPxHKnJeloyRILyvRF
PJ3X9Jr6BgasOJ+Ry7lBIc8RKtuptdzkzBUPs2ebMIv784RcKkMitKAuoHSb1h+u6ixx7sT4YvGI
ydc2Wu9iODuZUU1XwO3gXYmRw1hRTXg3rMD8lllW8NnKzolynV8QlkNV2FO/2B7KSsxr+x/kec0i
s/4SrCPhrOUakEoNgANhlu5EXSUNRbPSQMBW6bDLG7V8xAFyfou6MefDfd1pVxNnaIx5InyveK9t
yq7fpIScvSFE5dRL/7aq7T6yTc9/H0zfoM3S30gYKnlPp7vmBNRrNOWMQPD08ll2XLzswoy33MuL
7mtpSIt8kb7Lm1/erOMyZppPre15DTfIkedW1HOu0Kh+zt1HUk2DXe2RYgrYzWKhyRl8S/SnE9Wr
YNde0lmG9F21aUwarg8pKGwWVnf/ecZ3qD/rkCqXtyZgNI5V0nIPsIRHezOcAXGlHLmNb3+pLUm5
1XYIzIYYFn4igc1fHHTbGxtQw83bvZvH2T7xNxCzrWQcMrymC5DnPW+Q16YSvmeIneMlSaV9z7v5
aBXyUiB6aO5J4xck14uFEPEhL24jaVoEoEKNhPoy7/t9Ih82+L1Nutl4Y4YWQ/a/X99VhyKzAMYX
dCSNlQStosMD93IJa/4qQX79/dZVRujFYNlQ0VeaDD2U3xHdrxBPTtqlqem/qIoTTrBi5XC3obr7
QwqRE5rTBWuUYCuRnBB/dD1DLufC8TwZA9DywsR1TD/5GL+n8D3TqTVQrcf+BPjfYhEeldF4QL+v
my3HxedwPoX/TF7KgNdbXgXMgWa+YUdyFa6V733paElB3emm12zmuBRlzdUxtnTJP5cr8RV9pZSP
4e3p9+XU5ZfrOfMc2ttf4WJXuVjm3hRd++O27nlU1zCI69H8/UA5bn7gGaq89GXxr6pTsakbKl3i
JfJM45y5KTdbmHwvJLLrzwT1GbmIXz+Q9AU6HHodu9jixx4SaYxTNo8dXg6Gh8X2B8g9IjxRWm9h
SUjpzGIWLYri0294ZnAOyKxPPZadWMJa0KWJoUqUzZAgTMTHn4gFYUn7HpSoECwfelZzmtcGJJeZ
vHczYpslGA0ggrBUvgIg2du+AZgQ+Ti4Z9igWV/06JdunEXJC1hgn5B072QR85KtgdnNjNUy9FAA
cToO0G+CgulptMDRj0u736ILxkYssFTghMymjpUeGsRqauecIcj9QHGxeeeuVK+oHvrOc1WVVzA8
w84MVYGAILmBRu02XbIfbnHcUG02r3d44EZIsRN8steyXgwKWWuvPxikAlWY25hsmcrGFGtNBzLn
11svAq/8aJlMw9HfGF18/+//2ZJnyyFsfwWDMywJtIjElbrl6W+gpBbeKziAJLoq4B2yKQTr9cZa
3f9hU2kSou+LvoNm941nTOQtxPQNZcrCYhszORX/HoZFdpJXshh8VnBoPDBwE+QCR1JBD29Yb3pO
9aQ5kGBpo4OeHix8SWSRbpPZEiPD7CIANZSoBitgZcqvUqgjw/QxGrlHpWg5ZoXD4NJQMDWnHL7a
PS9EpRiffXUwbPplGmmn/88k5o4jlAQLOFkvHssdMsKPXIpvddLY1a/Xl6+NRWOYQwx1/HZg5NkQ
anZNsILji6aJtkGe7V+NIl4GTYp1ze6cPLz2sJRNfVqA3tbtu0KZF2to8UOIYVkvCdoX1i+DqYnd
gQyzKYZrg9rOmwutRQb7PG8/JSlM0Qj748qUqSI6vD3D+4ym2kb5UlXvK2SRrgIJjjBM4nWM6QyB
OfdcVvOAUIEskp7khaqE1VoDHtJZurnjmXU8nz3kfdvbuKX0D/cZGMwf5ICHqoH33p8fdhmPNIzy
x9+LIP6ZkBkErHrnj1qPG/aIdOMuREc+w0BmRfYYad97PxhJffEN32+0rDyaM56aj+T3Kclut1wD
2/2drktZs8rfTyG+TMbOILoPZe/qZnSIfLGSO1NjnSG28GnzhNkccgV19wQ9ghUEgAja2K5zN8GB
mYOqDVquTfvM+l7WQojpmBv8Ip3k32gzfFL8jWST7r0d2LKPc8tU9GLOXRAh1A0hNhfRKYBWgZa8
rqnGbi+xtaey4Qr4Y9VjcTHNpOIOoAcYrPRYUiMDr8abnnoBjnQNQWGUjZcSWSLFc1KRgKg0k9h4
eihDjV6M9qnlhEcN/dbVSu9tpBQnU6DP8su8UKOdp58x/qrKweP6vYydaBpth42bX2Ck0Mcz3mq6
EZdEp7JxhIjTC3oouHv/cNYcGpyYC0QFoQTvrKv+UH8liLeaIYW3GgBLB9Bhjz1llvlJBlXM/h7S
79vd/RSLpUPtkNI4EOMqctTxTOfQ1KvWNrZNHd8T/ce4LFW4D6DuD1MEMT7MLxpulN28ZAzItbKR
vj6Qa4Fce03dypzLhzvDaE7jsDfzkuOEP2ODv1sWpfDBJaJ2Ydkd5N804gnkNLau+4lHZSWeqPld
9vpAxZkf8JaSSAboTKlbLyK4AF2eUZMt2ary3FPGViX6o4feV9MGw59gJAQ6sw8ubGPsRS0MKZ1X
tgLjmt/rfq62cJnVxysksIhxRlpo49mPDTLP7pbhy6I8oYdUrNyPvL0vz3jwNJ7S7x6QIiAKw86j
Fwud9TZwxdVuQtMW8BWAvByjc5Fn7ynbxesFZDRI4hZWKgIxWgQHj/1E24fp7zA27QOiNXBb9Q/r
9OlIqpIMfjnKW1Ox0f9NxBJELhS/0nQzo1sp6BXMg7/Z1KWgpvWxgIVqbnE3dfJQ/9+JKnaK42Fe
vQt7cvUcS5AZiWcujFHVVC4hQQwaf6gXAH5X6FLk+wQApC4rBT/3YUy8+T4GkxslJ7NsjiV3nRGb
9hynNJ3QBx4vsLVv+Y7zBF0QJoc9RH6dWBmPA7XPPLbFzLblaDQOuIVg/6czUS5YAlk47y9V4k3U
CBulpB78ITqHVg/N3QcoSmNdLcljLIFHXQUVbVKirGTyVtMt6+CWkqj3MZ8C13TcmjWumzYZy2FS
wTSMi29pEpd1JU7cV704OE8fRELQI17my3iwhnk4EvRYOhYqU5TIFIjxk6jwqewGApEFJovqCsUD
X/LP+aF2Ka5ZLJtyj9a2ivY7WH4pD5F8TBs4Wnl8IprQGMSBmvDT9TpgrJG4LtcWAJ63f0Fu4mc0
mbntNDbBwiaSAkBHmhj2Twb9hrsVqhV8Hk2T0NVLhx0gAb0Vsn+TVtJzaiNqMVVyI5j+zdNwRNIc
9+Or5dPxSEILNfAQCTqZKUdTQPFofw5b7OgZQxeaJ8uqOQCPBmFnI90bukxnYK4DgY3k00dh1lYg
W/eq3RcFIIQZXdJfr42+Tx/xCfPEs+Zm8YnMuJ8q1ckJ71O84fRdweQjYfea3t68X6RHFQ8/CgIb
sn4NM4HKzgOptHq4hDwkZTO09/Q0QkOmWVQIS+2giPjQs6VJ9vTF6gLUKauTfm24aU43ZGhiD76+
3l0TTWNUA9XrPz1AJcXIZ2OUmfo+ICLuCiUvRj+A3Q2aI6TVvqucFDPE29vxZnoHXza2mabRxWB/
W+RLUuxowJFcDKlDoak2jgQ+QLSISv/DHu4yrmkI8V2oy2irY7Ch/p6aJZuq9aAU+iM0cFQRgNYb
YQdVUsyEW3oLEaA9ZgpHHrrCLvJWqpyqCLlWRf8tJY6JGPyZuBySatOhJtBHFwib3gWdGKrJVDIs
lMCAEhX2b/97OLKjpNPhy7nPXMUEmeU4nPKy8uEp4uwsm51sy23pTKASB6x2cpngLEYkslajmVER
pPWQmCEHBGHasuVoCzrIz8NmBfczglubzq9RkKmtbGvEBb1BYVqlaCf3RF2B4UKDew+SmhGcUCFM
mOKwKB/M/ioplYvbFK61VaP5YkgnauVuleOIXKeAcS4AILL4do0Poc5zfLQ7utf0SMJr/ni/zwMV
x2wcmpGZJ4DUcQ6pdHWLkScp5sT199YKE9w75jT5TnQJEjP9w4qJUSZL04qPstkJxLQMFPJrIhMj
8oS9iJ0iWpt3U7sk2R37B7xsQC4nUd8BXEwbqQaM7wHxD8F/zvJOuEEtE81YbzDPaGzFMpmfWg/g
YKxPofM3Bvbu99gbGyYnFcS8R/5XXyIucpo+KSzfL0LWMJz0GO84XJ3dLXn2vASAsXgQumhXYJOw
QLZr0QdqfbHhGi+JqWJoiBhuNKFyL49xGkrLLvNfVeiSmJ5ATagdDDPkgXc2TpG/Ys2v+OPo7KaA
faVk+8k/km22UTaV0LSPtGsYiTfz6UBn+2KZftLr6dhSwz/hGfYTqooS1R1kZOeYTyWFVK4NdsFo
MxwhHi1eDnm4RhanZA0PalHUcuvtn0x3OwTaLfImFb2i9m988W80yni4EkZXNI5rh1Zgsm+VLkva
0w5CDMr56/iRLD/IaAkLfVm5S38a/GmRXv4ZgnzvPrcUqWGEcrOZ+HL+b06/96QtxwHBVNnWgfjE
IKv/W5kJtd4GD536vah77frvq1zj7B2HE+Bs1tB+ANPHk150XDymiwyr5htRBtIoQZN4pMAfAOTR
hpmKy/bxUhAOl7zrhmke1uZZF//RrTAAe0P3O1M+0I+miCC7JisOlNs1nvToePZJEhLOxRuS5Ngp
SiyKWAHFhfARL9knd3G9hsq5uhlnm0AMT93ep+dyVeyjqXnrf2zqjDo7gGqDvNiZfczzelyBsHHS
HZuhRXBCeOcv9dLEumv/bi+3KSCt7T8Y28ZXFqG2BEQ/+BMyDltoz2Olik+0tuYx1Pk6F/2gZlZA
VumjBFzPqVjtJWHpb1Xoyuyz4R7dmiptvdyw56oeIt5AqaYbmZU9u5hdfnbl6ADTK3uA7OtoPwWp
QST6wyZiXOoaALzNhbCg2nb0sLkLZr+82y18r+VBbbmkNhG+Wyq/QMNGwbaopYfP/oTCfFzVuhDy
rCT+7YmphS4bKrrtSZVGu6Z+lskF+m1JcWrZ/B2VAL/6W8fuLUyxfTOlk7bXdxrUjQUaGhWcLPg/
CKj1xV5G4WiM6pPWYH18vnIjJMVxYRD62s1RTbjMNxLegMKXJZ1oxway4PRM+6yl55oUyceVlrTz
LgqJVm92veXqnzUEpNsrcbOtiHzsB1vYid51oNWuOPSuTeL/9UybwW8Fa/Y3VElXtjxSqCv8YbTG
br2+0jzHyWV2KmOSaxgDv3f9Cwno4iQRmAxC7f7xPau7mteTd+DfN87iRFwG7P2B1jq0QQsd22JV
U1LcxtPwEDOynv417QumHhkua+RyqglqsVXZtECBHSnRCElfKIG88k+BUntgI61Uj+yMlTYFd4x4
9kyDZOPThDqhPFqD7ppWKwOWVosUBTgY64FOJ/I+OGA3F807MB0fCHhyYlMQwZ+OSNuujLRVl2e8
vBCmK9+HYBMSSLG31Oenbzot1m2GWsJ+cLop4Dkwg7P80Ja/S+AiOXlrEVwodXLObafCnnsC6s8i
Rr/XM2892jpEHQYNQX+huLGghXrbxppcKgHJqTvVG3JVgkPzqGmO+P/xrz3tNp+qZzq+Z0XsZFG6
yi8ubaRxbk4T0NQf5KraZKRoyyC+hBLzvFgWxmgI6QU8cSf7bqIx8hZIPFzH4lzNfTvm3Gx02hx0
4G4Hl5S3ucTwY6S3Mr29tYZ6J3J9JDCeqF7W4r3SLfhVHmBDSy0O9wF/1Og4J9OmyM0/ptzniR31
pX86HlS4N23SNse0v9GJ2aSAd9cyzupJkcJgJwLTyfTPCU+PnWMXbf2kEIvK9TrUQuIHoGMXG7Nw
rPccIsuHgtw/ZfX6QAH93Ev3CO6t4cYfXnLEJzukynLRT3OsgQfUixhChDGLr6Wx6wFFEEamwCpI
Uu/HArcQon76hkm1kuN1yvGossT03zOfPNXi9LA8Dr3QOA7FvNMQNk6+PytK6gP5REwHN6D+Fv5v
zTqIpLJPXa5cCnIaXyrGEBnRxxzfP3LL3AHfU7BdME75LwVmEmY8xfpG5j4vWL7bxW3FuPGrm0x7
WcZS2M2gqZg4VABVShVBrhJHDMYEepSEoGDXuhNvujrD+crjgxmN0j22Ri3vSm4Zttb3B2pDaJst
5nDOoLkFJykzL9a/VJbPz+Vq33MIoDzyUv6P0/TuTF7dALG/0r2NcpyAe+Uz4E9F2Th6tDfVwVXr
fB0x2AaObj1m1t9rUTFNtTT597+q/q1BvuUQ9ToZfWHG59XHyBIJw7U64zuO1i40l6zE6qUThIMW
a9dhb9b/7D7Y8NNA1MQbdTqRYeMdKp9Bdy2pj6NPqMf3Ouf5FiMrkd7qQS7VooWPrEp6GH1OMhda
X0kI5iCQiCyfACIsWXDF1uQFA0JjIzFrvW5sTjF2zu0IBPo/eIk18+MN0j4XKHNgeKciKGV8f4UK
ejxdmw5CYZw2/g7zsMw18KgYX2Vn6xHiMAQarwNRatsoqhso7YsfGXZGKnnGKh2JFWBLSYcsTkJo
ZeDCwdR3dTQrlSBmIBM6MLttS5tmvwc2C32b6ZyQxmFSn2FnQuzUGhTRqWA2252vCOTOo6E4h6S5
DvUfbgxKFcBArqNnJ5xSFTQAQRNIxrzYz6ajas3u8pemOs91aAq5nR8+qi6zZ6pM/Wk4JG/2MyEm
y5jfwTrZnQWAvYKlpZXQiVm28gQ+oKh2D6nzU4ssbYCFkKNhd7EiKe/vOCd0/37oK374P/u5Cc7F
V0GthTM8QxjDFOxzR7WF2fgVJdN+9EKg5QMB1In7gIlHQeuRFsAk8FP1SNqsZgbkcFdirDCRB5iA
HIxmuXbIgX4BHJYl+XAgOsPTRwMCs/i7Yff4Oma39IbzXMphp8Epx3QdMVyWJ4KAvotoshHsU7xD
k8TmoB2IbaP47TxvtJXkgaWEV/kOy9hLxy35jP3IHNJ7iXmqjcMCo5+HqUEN/ozCjPPPk1FWazVr
vfFAJIz9B7VzwVoNS3357jTrpnttTcuDSQUlvNsegdnN03JSPLQceJzsRTaJcSnw/6i1EBcFX+Jj
Fe8NVjz4RSfgbtNEV4vxoR0OUf2Wc5XAmDJPDkZ0PilW3bOhFwIpjwS1EDrsDwueOW4Ls6U+1IZz
frZrTTqlcLDhacRlr1GVmqAe70L8zPhRJqhgJKkNibZQFPxhO8/GqDczTGTaOu/8LrHvAGHoE8kM
dFKAJTh8PMHfFismNmbNNHrj1/PlsE+677iLvXg4FLVxDiWIpC72E6PixWIH2TMicS5mV49k7bJU
W0wm83dCJsEHO9+tDsodbTdn50I+w/kKmBKlweur3bynZLxCvy9jihi/7yM+8cqLRnWcnBT2aUpP
4RopQjAt6iOFzzpnFCQ2FklnIXO9bIbwsqf2HuOflRoeV/djB3i/FGWz07EgvazAVQTPzc4gfnVy
HXvnlWIFTX1MkZV6evmAhkZW+aca/yMXHKlaaS3AEH9LvnpVx2shsGE3zXeP4whvX/9vPRdwxwce
xk6Z7vwtnxJ0WP6OybdgZ0OKSaXM9prtCwydKkhBqBh2sD16cU0kYZ/8FIiiTpI7f59LDQ4FKzoD
0sb0JdqqR6Mn0CHyE9IcPoDaq5LO/4G8DKoM5k2uXAU8orKtVxKdvcyTzyu79p7EsHiwW1k8c06D
RikWKZCgLH04HVvZRhaDvyHZCFCPRA07Ic7QsBB1EMKWy5sIUi8qc8RiT90uBKUuEdacsuo3ats5
NHdRfoDjnqqENeg8fq1Xbba3qIwertGGJGEL2iYc0V2EkxD3jJHqQPhad7bqsX5+7a64OFCEFcCu
sdBNMtX9fHqCPAAV1ZIKqHRMTkBO5OJO9Ui3ckJWd+ttvtMU7IZ1qmEM8vlLYEG8r309jKLztF6G
0Yqi74cNW+vkn0JFPRxu3bS8ue9iUElv0QouvCDIekWbtyYBtNZ/OpLBwjOR5ylN0jzB2FvAOGo6
NAbkgcSNMuFZIYOFsN+nj0gy1hr5x7GiALRTdprte/yeCiW2VL/Tryo4cdN/gQUr9OnsZgQQchMs
iCXGrpJ/JoXqwPIugE3TMVMtjrus2LZ5U0SATQtbDjcLHMp/QmHHephd6DUuqhd6EMKQT1pZGjZr
G95FH9im3Rpm/NLpnHh2Eg3Tynac4T3jlnjZSXQbGXDRTadqTs8Y8H644ouBQjlO9t3CNNvOUQVX
ti/DLYFJsfeaNgVucJRejLgG+qDRqG0pOtf03bypZZDiA5GHBgn1JmpdqTlTW5D1VUEl6bnid4sX
tTWcmUCuKN/IwoLh5wMLp0gCZOXtK6hfJHhyEEL0exQ+PBdw4Ft9IlFX43biF7RCRrSKdzky7K6s
p2OPE/cMDo25NhIZ+RB6OkrZtRjEXgcRrCBeP2vFcNTjG+2eAwADZfZf+Y1zlEHcMH3B7Hhq7A0m
ZzK20uAPlzHa3LqC5nfQ5GKCXIaxu2TBP4jLi+nUERNepM6r3mwUHX4bynPaZCemyxBEtw4j6b4m
aNc8XU7ME44fxOBLNxGmFAMkxwQ3B/QprQ9fJ2TMhRoHkYhWoJmeOk1k3JuTsyJmZmTdL7Ig3Zig
BkcCjWYIXlatKfuvxUx/wJ+JMb0HZqh1Cxl5ZQwXPIXGfE+sZP8h4IQiI1r/8qSSZNlcd9d5Oz0z
r3v8G7t5wvQxRrPW3GddakP9kchL2DLONwdndweBSgpg4/FqvMGsnMy1I2pxymPxFQBuEj2XlA7c
XWhIyZdeJau2+AVfRUadPZoosNMNRPtOHsQV2Fp1t1q4Clqb0Db9RiviwikUYn3h2u2m0as2tXlw
fv2KndSQeSWUZl33ypjIruBh6iIB4xaj7USIVOWkiAfoUEt5eK5QC4saq99w95FChbCjskibyQtI
s1hosJRO+SXXZVC/Q+3k2whZj2GCE2DFWQhvJX8hMoqi4Qxzgu314P1i4HujPstlw3GSbpB5m9HW
MgzMUwY2ArA0Ua0V5HfJ/m4TZg1b7jPi1O539c5R220AMAxUF+3iZAcdHOQKyPN843z86BYHpkM0
nLsW6+lgXoFUWUzFmEVuPVC3vnv36IaUlyeUW7Y6P9/D4moq8dFKq32vHfXsjS6mcK4JCghDycOX
8hbx/VvlEgO71g24FjbOEi12/Eb/i92IMYCNdGRjDnLypxjhsQX8Dj1op6Vm7nfRjinYSfByLzdb
M5s/eO2rIEoXjZexklGNyKSrRwWAckuCQj7injHuNJ0zSdSiWibn83wnthQNwQvKJS74gAc3mna0
VWi9KnfFdpG9RYCm3si26YEY6GJO/NrZMlRAQeDGaqeRntl8unJbzdmo7W0Eu4d5b9QGrltAysy+
Tg2H+5I5Q6xNomF1Y2axuENAGCJjm2VOdf7np0d3Ya6VIxs9Wnnie0t0FVg+W3jfHd8ME4IMn5F+
c/Jsc0MHN1tAkwAk6CoxpWzqhyM/UgfZmHD2CcqU2XdAG7kbd9VhEC9ENrX5tGR55jGxipyilq8+
O993QfmQkFNPGXehgptObQ/m5qjDa0DU9KPzqASV35DN9sX7/0XviOS1Xs11WhCOmGK8M7ZnQhw4
2lTza6p7JegooPjWxH2VfeQ7vfbsaGlalY/Nyb509/EYO/xUpHp26FkucGUOy8xGDpR9p+zJkoMj
twQhM4290K53z8DpbAhfajpLdPhOUHaYjthaR7PkE7W0+BWbrpixdj+asXEGhHdlMtdyFOvmMZPy
qq6ryyQGZKNRleAbcDoOAwCvorQ0wFt64qtg6AA5RKW/85vjx7yH+RYxJxSddtAfFrWq6BG6sb6n
BUJGvrw8sbQiI+B0ZgRm5XxZabmI7lk5lqrU6y4V+fMNAS5EXdEuMWPgesu40ZV+ounjLU65K7oc
sW/7TLwFTB1UFATnZEu93yAVsijPRbyjIIbENi8gH25c/2Urz2+pCyZlRURT73GrYNNSQMktmRfm
kjJi4mMrxYimtyTjp1p0FzexyrvdJ+jAS5jTeWiFeDkLy3hDCg6T2r2bZLy0oa8hnn7Ine7OHfWE
HzLsUtKlk5p+lLgrLaGP/u3YQtYgsXNPMFOJZD5rKZv/rZMwz+A1uXVkSE9c3GcTftsH4yUCkTvP
fwwatBFy2srPsBEtHGmdoZaYQesc1ON94k3E61HK3kWGrZikE7FEqgOGQEHi4pyAZX/9OkPLkrNV
SH2HIx4hCYtSyw/vhow9CLbJhKGrGUgjTN3jWX+S3zYzyylQUFAZFORwOxaAlXLZhTTi3FMItfU4
Zxqizbu0nxKS0PEyKzs/RvuOZ42Sh8JPBrLeDB4qONNFScKhgZWH7h6REeTGIAjjJ0DgCQ5QLpRi
EIs37MgaiRqECikZ0Qd5pKl03E5dBcuIDsOj0MR1WAa/u7wUFcJsxdIbiIRVxcT84xl/gEE05IY+
l0a1UY0t5r8+StupDkZzvnU8SFn7WZREUPrUDXgw85h25A/Ifv+R+pqJZ3Cn2Iuc0wGnhEArAWSp
wL580pJuXNwnJ5cCepC9uUGkP4drj3alb3vvJkd1xbeCtX1zjkMptY9z6eM8RnAplk0quUOucbmW
VRtpGzCOi0wjc3wJoeyI3cpm/WVwrQ/ZfFz3gkHw2HQSaMl7xMKADI3yay0rFsQP4QMb12KA6UVI
Q8kWbqgck5seTDUT1tz+yyZ6wG1KuRsQLYSCIqZTrdZhABBELMSDj8givY+pw4iNM8ocPgl3lHz0
Fyeom4OC2L1zU9v+bvGJV7D4hPUcjgq3JsfvN2ctMEeghGt9UY+kmZTFPuQSfaRAeYZGU1MjdPBG
2fSv21lLTXRLupBMqD4WfH65pMstwRCzwf9ChrCLMbYQuO1GKNueaoAeAZTobWtGTUI8d7AIQh0C
4k5ONQEPTS6Ayp2FGXUD/wxzdLkw8hQ0ZQzLm4IY1UwfayRCp06Gaf0lSsF2lZkVehOv6m8CJZU8
1PG/EHFqNV0+QMyO9S9cj0zP/Hquthy4SyvkF+SD0Rbp7gfrNT6Os/V9nrQ9mme/cJsR6cVWkKf0
/7cIA0LVwznh/IKWhxa5xk4ZJLJKylkIJSfuL3yW3pDFOo3cjdgcHPKBOPvjNU7WbGboPruBqSzI
1GyHAiNMoQPOiqbszYo3lTjHaJBLddJZqtM3p9eQVXPU+PJn2YTWqllL9SwyY4k9WNUinyCsg6qw
RdHstZtD7sKUFxt0P119f7fRjOQOOORFLQapzYKuk2h730/fMTMTpg03fq0dH1C7FBcdLXLU5nuw
0VemltOGkePibvCZ5+H/05HXtldd5YZLAUF1eKeis77jHygkgtdL0zEkXN6ZrpkC1IlGZB13WUJ5
rPdyfQxvRrJq7X+eOVDJJeaJV8qV7cq3OXY1Iujw9fdW5ybpHp6aCEAVrOL+zB4wGUNr5YFfHlUr
TgI0jpPi0GaMv+au4d2p/qpfe/XbY6Bw1re7VXWClImqCHeT0DxR7ZzF2WMyzylP69/UFdHdMf3A
YcsaI20euy+P0dmeasNKSTe6+yqkKw5iYCwrH3Lp/a3JuX506XQmDvACW2rkzyXuk9oliEIwAOAV
nZtgH4JwXwZJ/v+IdShh3UXPS9eCoIBCyM/Il7QWjyomWt+50/cVnFlvoNdmMW5u9mosTofK/fkd
kafHnTIs2zhjnUfLxBwj2L299zByiq/z7TWB2InJ3vS0fW3AqReunGxMeWzgPbqNaBr9TLVUlyyd
B3GfaVN+lKEffRPnPIddIT0nEUdr9xM30khbS0C0iTKuPqTtOM8Xh+MRSGHqNT6iqDmC5eXRIjDp
8e0q3lGX7r/LwTtpKBsQCnCJbAIlpgfJQ6eNptaK8J3LdiNWMp5fz4iWPAXzyrALG89FOULu1h/Z
ciSCR7e3qSUmjjc31VG2ChEKW2XkC6ZcDIBPSmPyo+o+fIkUot8ETw9SX/x4+3oJzUPoXuzJSOWJ
E+o4f2Jm83HmX+8lVp+kISAG6j7dsg2F8boPlioY46iho+xQbumTjLKJN6R57BEtEX45m7or+wmY
xAA48g9dF84Ah7bm3YLNPf5NJPKUQ8xCKDvxh0X2l3pgME22ut3GALRWBPwLoMa0pom9xIpqY3ni
T5nPC+Pj91Baq7v2qTB3+HdFfFjJpYSZnfH2x6HWL7i0TTbZTIZ2O4W3SR3BHZ4Wyvx0FVRl28LO
ClgOWIT4GHPkiXVmLSjH+iN0ieNIBwH6UtcDEgrjnsJPcgsWi24+KH07nNeUQvxge0u09Rv+98vB
ZMKZ/aGsp740KloY/rh0VTqP4QfjB/2gwn3JK3Jmy702Rw9OJCvp8QlxFJrwaxctStQKn7UXaVRM
AUtWVaqcITNBhCWsV9F+7aKu87nMTrsRCez0ZmgwGTtyjEsCyq1PMcfsakeCCw/Ye8Aa1lX6rVRn
7XyMU+49q5xnQi/RDwM+5v47CRwSDl9QqEn1GF055NJQNxbTzHb8lx7YX+cgWqMSUPq77sn021Gv
dVLoDtMz5sAPVp7BsCdMyP0je0lb5WZxCpEeFtBA4CFuhE3nRebQ412KNsXHvRZ7afBb49JYSpDS
3vqnCJ+n0OUt8VV56iB4T2h7ZVLvs0Z/LzHLzeWjq0k2zd0DZt2eg+tsHZZCghpdn2veeaXdwcbf
ATsOQSFDj2C22IHc8vaxGue03XQFqD9BgxoAQ1xOs+ZlCGMglCia8bx//0DnbqEMw/QEcOMoy97e
6NPXljA9rnNMXaHYRIpYCbdjskFN4HvsJMl3tsi+bBNbgWmq/sw8E5KoIReESnX0pUBI0ci2wRmR
uzo6fXsh+kq8Fh20ooATsHa5qlMjNM26hyf7I6zGU2POfLSC8RJ1kbbVMExSVJ2ZQAfhmxrc7ZoR
J0xV9nlhczrjUvih/dE/JcPnYqNjv7k/HFnRi3e4EhB8HvUkMlRv+0/xXemT/8+z38bPRNPG3y0n
/XeE4ZiAjZlN3uLUVbkSHx1G1uNwzE9SvtlpCMzZWeCYuJkFZc5zM6eGSdF4a1+XLH9kcqULWf0p
zzhM7/dOoaoJsg49JKQ6o9vdbM7d3VRIvgR4GEcEswtyYprM+J2+e3bAAdVEqFzyX+Iza5y4TQdm
8tejMnEy81l7JplYIhEu1yviHBsmzkHrjCIDugtqT0exaF3IhkFJV/FKcbJQfVPPd1Om3l78jxvz
bDkn+CDNsfVJzeQ2CI1D/yrSPKTlyutHMfzZQvoGjt8BRb7RzFd47MA1SDkqJKV35JyQkWD25Blr
pB2Y3JX8eGjpYP9NFlekAId1cZUDV1WrxvHyGWS/PYtP39VK1lfAk8TeKqJWvb+jUCsRtC6jxdvE
6DRJAnpC7mBliF2OVwJbfPpK+eE45gLGr+gXP63D7MyZyi/KE2StPIbX4PxqWH7rxiFuOZrSwd1h
4V7VUEHSNnqWOltEirKj9DkjAC3tsPLOAkhO4wkY+q/my9Pmfax/+ysvEc8KuzA4yDjo2nX94mx+
5UgNwoPGPCCS5a7f2k4tgYc76vBl1npQjFqOmAAaiNGoP/84s3vgo8Yg/YbLfiiMkhiEBLBe+IPi
AvnEKXWDCsdx+HEazPC69w+CHxeYe1jmAA1jsir4x2U8+Hjn2LagqZ6OGI0u0Y3QLHICkwMdbc0U
POOkDfaHP+qd+wvQgntmlY1/paCmlCm/HOkhMpK6hdlvXogBoqL//1CCHoI3kXt7BM7mhmGt1AMc
or7+wx5xJllwZXEoYnliNAbN8PKHjilqPd+E5tZXfDw4H2JTVX0sQB0yhxsMSj6+YGxXGdeWR7eQ
lKEyC9oerKd/dvxfrZu2KRvitBOCOw4Vzg5fsAXYTLqejIwy0RAkput/xeWzH3yOEWas9Dkf14wF
9gZbMcqDaJiFvtQpmRog1N7XwgCnhutqRfkYAh8rXuyMF8jZOnITrN8+wj4APb3q+NEF0mSQMGlm
rwY8lf+tObeCNLVFGBUwT2J1F9dAwpdcycCxa0rWgEIucm0e3arlwgX/7cH7ULT3zxpflxi34qw1
Ij1qPM58Ow2ANYt4cZ8L510z5DjVJqEoHUx6+3OdptP47PlEj+DM8Ia1DZG6sfDBz4BYZz0PGqUi
YKnsCNs9r5uJSLTRZWiFooYFW7x0R5bCluCtSlAZC0UKksJJqvmNRtTIIO4KR0Y1A3eONtVZUhcZ
5p4eWgIQqqJYeaApAA/ErSuPyYWdPYK0tXO3Q0QU9LZ+YPH7aqyDof7XSALKpFlE+d7MNI8MZxwN
rNCmOsUHfiTlPQpj9Hx/gHddu1afbJ8TAGHOUBYYWD+tKti/laDiTK8yTAJf4rC4ULSBEUp+h6Xm
IUR8knKdnq8W662h8UdIE2efOcWRK/RxJVfe5VsjT5oagJfWW3T7MuI+ca+Yrzxn/npyvU+EgmAT
9+dpxYJCfVIBsPeKt8W+ZHWoNGIV6Ewlq9+1zNbjhXZNqux2zuDJfsHXS6h22eKNqHQvqwmGNBpq
HCTSEm2DeOzHyzebkPGauP1GDQFxl5qo+gOTV1OVB6R741zoKLQnqOdVV844VyL8lpM99uq5QsOQ
Nkao+v+3jMaLsJ/dPq6g0iv2INgOo8Mcj7yRlSnWp/BhC8/fztV9DsmH/YEz9tP/xl58WEbjq7i2
Pq7GEeWPZ9/JXdRfN+U6r3FXaK0hh+WtdXXb+M8IvsDjld2Amy9cYj5GQS/sxCRHxEHzWdLSx0SX
rQ/4hiIFXajtc30pI6dg6Ly7UmlsS076NHzoK4Bro7V3vzj+ygGBNQBGONuDNhdViV1KjPcdRQCN
etdm8O9ORGtAGdrz5dYQGvAt3qC47lITdFKheJvVTdTn8SjC4A5F8NYDfKZ1ZXr5/haOx3i5DgbC
G+lAhE7MhcAiqBrXPCORKLm3x4A64aIfAx6JfZ3qiNUlInM6iaOtro0PPEeXGwVrHWPsZgII5z5M
tXx2FidM6PYAesMO7+prwajDv3I4nsdJ38mQjteYlu0m6SQWwAQ7dR2CRfu5qAd1He8nvoBLGK1T
c1VYcdmbXD09kY3rlI2GzuJQQLnc798LMzmgWSMSCGrF+NT/tmLznkOrrINoBYM0F7IWS4fb8XLC
iTnmFo5a/yMzc8748Kl0wENzP+n4mk9BMXf3NlHSwDqPCmUUNh5nFX/Zwk1FA9XtyKsZxj4wn3VM
lrXcntkF9rOm0SFf6kK/38ICYLwr5NY610BdoiYc69iIXaMyOLIiCbdnxYCcHiFiWYURLvZGMmff
JcMOhmCVAto+RnbHC/5+cyXPuXX3KViUubLCdvkReLgq1iMgAzEi5PiUnDfaUkGkY44JVZL6NsXy
8sNfmqS/VUJHkbBNle8IJPDMVMCC3Sj3bDtZXFCHT9jIOARgPfOyR/3HTHJEqzc+RSZFzT4GVOjf
66q75MndkNixSLiQccsTyq26JulRkFrC+ki2b0+UWU5ms5NjNHKBMtm03UzO7ursuGC1MCnhgHrX
J+eaRFQ/q9+RLsnNePIvd3gEBnVmrrkSLxAF+wBtoOqbTZ8WZnScZiFNvPe4HuWrQkmRm1Vn0Nhb
YWzY7Lx7nfmNn+dvweneokNH+M9APHhosTHB9BC2mMwajLmpUJaGCMbIDQA+0JEwG0lO6GPcrPnj
9mri3m+FiGgNep+mJf7Cg4kkoqvb7wFACiCTAF2E0B3mJdUolI9b/7VThIEc2fyrrRaYYy6e+2gc
vml7tfrlBffKDfpkSzty+ASQA7rp/GMlZ7UE+q7vLLGtd+f12SnFOrnVxuHSKRh4cRnStYQOXv4Z
oTC61cR5vv4MPDvCllMamI+eVD7Dl0CC9bwCPY7jYpJtdUlqJkZRM9EmFeWm+vEoc4bm+LnIF6ck
SY0RPqoMmqBJHTNBZGq+DtXVtuykX/xS0EuaBvcxpIqA323iNz9vKS8MwOepW+8UXBYZNBRIT1K9
lAt3M4tCelPUe4yILCbj6RSSvfOvqZYmvm67TK9c0d4whvOwy8G1xP1h2UAyRSj0pXLqpMkU3Gik
Gaa7hsHKmKk2iELsFAJjn1OAWWMn1QH70cpzde+ZIlTup4peQxy3GMsuqbVD/v2T1g7YR4DHSiPy
kJm1mMx4OoM9wTzj56ZIMGdCtGtqvOXsa4y97VRiAgg5nA40nsNobMUHQpRMH4/ILzWiErAQYXQ0
gCu/SEpCkILEMjFDKGWnrDF1UL5ANTiEQIqnD6/k8YkUBo8u1XTLCIapoTnoK1SISOxCCRXz3bKY
WwFzeO/B9jeakQAG0l6bsZUb6REyxdcnq83ATQ/RLoFiF/N6FUrNNLfP8pqxeIQL7wOEXlKE+jNv
oN/HypIjxESF/ePX7n4yApIy99NRVqCQk8GapkacAHIadcJfLkRiajyCyeUcXSVStVQ27BcnK7OG
o+IZqCDYe2lDQ5XsVQnpS1vkl1gFAFm30EccIUKflki2OLcpoDpc/+6mn1fsmov2xkwdskW5JKqe
kJwbALbYk7jEdKpwwa/EicVVyQxEOX1/F+DJous5GwB76aQrW0r7kH4o84FNp10pM02FkcMWXijZ
w+2wHqFg+0BIxn23FkYaDE27ZP3nQuKfftkQG7n/RZGcONlevp2XaGFyv/j3+HF0OF+2BM1riS7V
zngu+STGX+sYFMUDqQJOhAL2rDVZb8Pms9gMf9DAYeds/kjBnaLnNB88Vuk/JGuubaPOCJC/8Xea
yPtRUiNoRYc6Sm4+WZmRPlpMSVlwelauA45UoDU+5OLHpKbfECKYRN9aFftEXGyALXErIzW9dRlP
3yDbJCBiN7bh/GLWl2BM6DVqIcdGPdVeh0ZiTfyFBZzbwN5kVYDHS6TMhGhR+YYfCvnN5WdpIXLA
B+C1DSI+5qKFEE4HDN4hjiynCGnfmIsN3fy49tWZLWHNRO9y3E3POu6PbF8G/VJkGXzdV7bTJ0Zq
Z0g+t0F+7+n9csddc7fgk6PR4Hh2tP3K6stSuBN9EuNMq/+5DMrJyfs/JXv2UsXwokEI8RrOvuVL
cV8xrRi86RcCT4Ki2lDubZgDI4ubUzzVvU19+BExgle8NnyK+6MnCASXLY1ycBsz4yDxQQ320U7/
wHFw7R9GvVlIpNjTOys8SMpNyVCUFazFqka4dvzCqPVaKNhJqUZhLZ3+QTvqbas/6IqAHCuOeH72
X9vvNHCOFmX1Xh1NtK2yw4gecjX+p4sb9q7jhEbHeAMwn8t3Vz0V0TnWpdzfMhCuJjlcn6y6lK7w
hRtv3DXqHx+J9KSfNULkvPXvpEy3MSaVwc0Rs5/Q4XDOX+1W3UmaOUa10XcYEALcXhQE998Wuetw
0M00QBFDc6thfZDX6pvdfVrMrXjuic9Cvfuhp9UykGjPWODq2DNpGTJ+W1umXwDh3ufernr/g5rf
ck3prej6noj3svE/E7kxFtzcOwxamvDfIqIgw4y/VIPRdIvPhMvn+oub2bjkCgrzk8ro6ir8gvIV
4tYzAIWEpHtuqsFi8/xcagf28kmbBdq8nBUpUdNWLCwkv/JQqFe/otTzX5+EOJyXs4j/k0HMCFXt
4w7+AXs+L46zu7E547IyJU6bq8s1pnop9MDKKZ5hH/HF0NQq1NmImz7MukvLom26+9KQnP4bcWV6
48lsaMPcVx/byXi/pTCdwYHKP/SkNA+0ZDTVe+EKdXV3IS5FBAz7N8rEAWcINIxk+zcymJWTOdUi
2REaPlkVp5tVscTZdxQ1zyIKMRdKQS2O/qlimapHaN/VSc98ns3TXHdFvStUGoF4bPQuEIoPWGQ3
WprURcmCO+a8h8LFvCabnMiIR/Yi2r+/rXypi9/e9jc9YZ8yxLX9hfNq121i8bDeU2lUNLIO7NQd
A+FeNMQfDmFPBfSggf+j/oB8mPhwTEZZ12fpxcyF8gyz2DQk0cbhAoOH39CjHRQPvsTscVhWM2BR
ViS3l4mqaWDSQk24mA6jlQs1S/8li0YBhnheHwlaBlUIcUOF1ajq9TiX8A/vptBp0EZX5GR1w0DC
e8uCO3HwVfYtUyQO3z0XmbUnwhFrZE77d7suolakDzktr5nlzbqIzKMPMQwgTFaN4QPRGzd+l17f
18iq3Gw1WIJWOxQAzIHqDRvWSGy6wx73TuMXXGxS4XHe65EeMCh8VAlpVcHfg7s0wXbRAFhhqzaV
Sf0qPOOdxWDMZ/qBkEsBA/atCPagQHI2+9nRbt+MzNizAIFZbIgr33IGbsDf2I75rJ2Sjyn/wKwa
X7ZLLTDDUxPFtRE5/WoMfq9c+otV8nkfs/2EDwpqwxYVc9QyVA21phLhn7nwFi/MfWq+M8GTjgY4
sYy4GzHOGgcoZ6MWQwYAR9BM2x6IwGsXJ5/IWrwBtkvq9HK0BzgOYQFJNHoWBiBUvPcAx776rsGh
BX+l4x7WDzuGJRfu+wzDxjS3yeqEUxXzKJGADVXZVT4/hdSKQWGSW2lSuWrX/+8aYH4xD9Q7ETxf
842+sAMM+6oZlChC+GaX9p9AMyszN9D41yw2iNEImQ5+1BaUelELGq7kbASvVrRiq4khBBxeDIFg
bqNCQBb15uTFJXH34FBgGOLhpYMRJpSOVD2oc+/xaDLlTNveXSKLp/dnlA4PfYVpv+7bNRb+Hue0
Ar8kq2YJTs9nQj5WUeLSKq4PT2ZcyxwaS5av0PNXPIkoWnkcIY2ALCg9bL+Or3cF6zNkj4kUxoxZ
En1T43dkY9PVP2n5IyhXduCpqY1s/mKpJDsE5ELx+zkzVUQpb3r5jOI4Mpw8/3Sj0IGa7JHXk85H
DtFISMuMMSxYkqn+ZadPNzft3WQWE8Y1uiSFYdFAXgk5d5ql6HGmJUJKjnMgkGGiTWaHnWADw0WS
uplvQY06Q3DZWSzE2NOJMQ4i0yKgtmiq49iLQjrU1eArt3R0QkfZNy5gWpFc8/8QHGzjgWkyLS8n
rw/Kgik1bh/55YfhygVsZv4DG1y13EKyZYNzRjI0hQQC4Z99yzjaXa81J4ncagQy7I5kUHzavbGY
9hoqsy4dDU7dI2nKFk4JDzNh62mkgaLEemNP4hhY713+3C14+BJSeJ/puMudrF9EH4cPVDfwecPS
61pOqYoJXpOsKm7CHWSuQwZbznvBGBhrzIfIBCI2fGs1oacmXu2Sho8lksDsOoih6kce5xYY6lXr
8RDPUxJYBMTb3WXr2lfByWcE6UoCd2n73K1usckjLK8M9ldz5Wi4lWO36V98hqMq/0He/E9R7rAJ
yhLtIIc8tEwkELpq8pizi9+ZZwnw8CDUnFXoNRhWBfdzQE00sswt67Pdz0c35ZmBaY1/tg37euQ5
zHu5HL1PYXTTknzWric9vhIqYk9nPLAlDkZzSNt2ghap0gI24ZVKD1ncVgcwSULV2iWvd3FfmZ7T
YrOXiSRuyE9SBjTusXEjvBfVZME2mh+NJqvNSdBCDUCOgxoEZrn0fRMXfBzcmy2LnPRfPJT8g66v
ZpuP8O8K9PTLAFfuEvrdgtVH4PHTNN+isw9dOizstX3EtbqG06QehAGVr0EpkE2awol4CN8UhwEg
lVtVAx4tBsApwqPmo/eLaZ0zLkuA25Jh+po4BnL6RSEnt9634Ida/YlJ5CHarSvxNUZEKWVC5OFH
W20+2tO203bWQnLVd7suAD4DR3/3IPemVpRQ2X48LVXRZExwIpKNfYBbxaOU5yKn2E+J2pn3dFRB
O9fSMvuNEzNul8fIgODFgnIsKvKp8baVw+soY8I6TQM3YqV5jSxcHacCT5RHePNs7uwYjHxsfbCg
GM3K2I58oXV2vHOzSK+sa6xJAVm5xT2UVP/Es2us8h3vkdg5A4uEMKop5GWDhQszJL4o+D7/Hy15
fA7HgfUlZrvXgGBQZipsYSsjSrSmkqsp/1KkKdgq4QFkFrwxWc4hgbBw4wCQVwrqTBvKNELKVI4T
F+iJ/5KZGkdjYYkVQm5Z2bm9J/Z3XvehxeqStEmzDcPxly8wTadwLPKybpOcI75jwREIc9nV1IF6
wvd6OVyIyZFLgNC3E1Br+US5wZWXIuMcYGaptyh2qmRYc3oRMHzNe4rlEcY1btRD47yFW58dOAle
TJbOenZVNB7y8sesyxLrQGPRNXbwYw3Nvfn+XI+qrdJ1gOoRN9RoHgwDWlXmq1jF1isLcXPpuK+i
P2WC9sD/0bILM3f1Z+850hmHvijnhMsKrw/XnU9ccok9BqStUO1G5DGF0VF8DsfBSWJe6pE5gwg2
WgH6DW5kxBG7DddmVyaT+i+TOAhIQlE4lEjB7azke3aM+Wpe0Tz5OLOomUs5TVd3zo5XoJauE0Iu
HtQw1pnP+BbUCGnjkAsFIXVgcklkJ4m9P6iPhU64bPmfYAhnwy6JxeCJrfxWMy1/CzMuwFv7YZg8
Ips2LqSq0nGuxff1VVquwAlToys3qhOkuDaM+maWB4p5KCLQuAD+jawwIyiNR0qT64aPP2+F8HRf
wRIRkzty7Kzu1kp9M+rOHqxhluWRL59xLWjjMi8i6HIWemHbnQ2btGUpKZjgfWlrtI/felS7LyTS
8LHZQ9qf54Mt7mSC0ZeJY3fkGg3kQPpvfHKbNrdjBu2ooudH4vqmfvZ/EtdQPedMCEEZjlYGhlqC
B5IS9G4anlc3MHaEdoSdyOcb18fWovSzMxAviPoOs207yzQvFodWjViCDjtwMEBlyIy3GAsx2m/a
tpAx2Waq7KzBPWMqCzeqiw0XfrTh0ujpDJzvBvsafOnJhVoVa7eCb7Lg0mFJbNJcNJ3hBFu1GPDU
vBN49WqgO/MPQxbM7SIt1kvSDiFIwmal3jqypDcdVo6yV57KZPlwJSZUD/NqcDX93XfuJT6iU4Kp
p4NYdRv+1mIQxqJxsMlC7jZ//Ps8aZbw3bW9aJjMbvZ42trCgQMU8YRs/14Fz1VCx1DT6yJTaW76
ju+WCqAzg6eMIi9iHnlRexAgB+wC5Kc4cRNok8aP+XHA4aIvQKruOwr9599CWZO7IAzfalZMnPrZ
V8IUvJ9+wsxukqCPyn1JNbbsgZ2KSjcwps7dWYwPb4nJLITsVTm47VhrIm/tMg/V7ELmcI4RyaGF
3A7DsT1OgSUXWZWOjOGbxmbXAIc8zJnmHK4b8E3o4I7IhV0Dz/bhtXWQhlqWcHWMKK4OaMY5DeXL
B3GDjXCrP6LBrvubFkINC+iDWhEkRqrr1O1BaVfOjRWLF5QXSmpUi3Oul/3ogI04SrdAwkI9AHXL
fjizZERjWDccLBKw/H3/5ly7Toc8cNKLJLVNbKKwo9nv1HU+UwTrzCO0bQ2YJJaah1cWWLNIAIvM
tqSKjFNXP8ijpNtoaJQSEoTVgl9D4lRkh2oH/k24/NwtNDdwvb+/3va5DcI+feW6mMc0kiUF3qUv
L8NTxzFlThRAUksKWSfanywQ5ptIgfY9uFyy6RJsz3d3TQikz6I7Ji/nl9l5c5LQ9vC2wxlvI14e
Ho7m5LODoZ4KUgv8ppHImknpgq9nMAQWVfvZSXSPijmrv3c3p4ySTmc29asAFvpEMphwxtlPbCrI
J3dSj7e+WaRHiZ5UED8nXvKC9Ccl7hlG1oUBfw7ZhBAjT2sbV+s4kLS6bfKUGfmDWRTscCRg4LGg
71gR9FD2vVrrkK+JViCZNkczod7VYTAZwYWRBuymX+qLnebywSLu7MX9iWxJPQs80i9CIwxr8B+x
4tjmevoFolN7jsUMOlvoE5jrpWfdr/NTGGbioI0y+goSZ5hdmEauMTUDoi6HdU3ljcUxNEFPqmAg
79m4JMru5i9LncJXjyiRZzXAI9fhEATdI7WEQbu79VJyul5slhhSZZuzKExn5ao9c0NdfxjkqMbE
HKr7Gi2JBx7wVIkFwK+FG+dP9JA6FQCiLkISPedOovwUaXPzxPhA9PYBTBPkEwAO/boQInFqQ6lN
xpRNfvngzEOmRb+BZJrYSShVBsHbbFq7+LWpHpvobZ+ACW1gEQS1PzFFXOTK7A6iZGj9MFjPfagb
BqM7mYMlAKtaHqZiPuZ8wmml4LZGUNjiUV+xT/ETizkG3oMvoIy/kaNzyCd7jbYh5A/Gbd66pacj
RQsdzZI4iTmhWHv14iz99/1tbkNzwVPsfgkQ7zEvltnKaHVDyTfdVJvMhXkNKWagLBlWpDJkVrZy
STK3JaZubEzfxHd2oXJ3aqB9YyYkRhS1m9CuxsVNDnNvxseK9KR0KpsiiER/7aQzSIhXYGDLVkV7
/tzyMRQCfVxGzmLJIHHd23cyZlheVqODh57akyEjmcTiozgco71koy6Miiub8ymM7QVZP+VxKfqR
mWjjDl3icitouSB9oWLjpgBlN81EwbgIN8OfAcanA4ujy0fu+L6kHKmc4Qx768t7fNiEPwM3rmj1
bQRVmcJm8+71hLyTv5ry3ARoevStQbwY46kuPf3qI0nnj5lg7XZL1lee9wWhTzfIimY7xWLRWxn0
Zh8FiW9nWhhJsWdmqttqJwqBXBqX+1bPh6sMLQKc3rcgXrRZl+KlnxjLoXeolkqUfCBeYPsd343D
kf9F5iFFfgDWMRwmI2oPnOmWYainkQiW6FGnKlYtdBHzMuegsoxeRW8yk3r8XO2T5pHfVVDR9Owc
Nz7HMLC6/B9N2eUCLQm8zs0ZlMz2LdI8NPPOJp5nCSnoYlJCdh8RwcAsfy1LXsDMeY4r5D+3o/gZ
Bt/c0zn64lMUzGTGKzLvUPcU7nQr37v4Pl4k9Bki3wOq+wSsjlBCfJH6w9REgPPfbzzMGviUD7UG
D5yvaVEakPs5K53eTAQ+Pwhp3E4ejSjaQKx6ZHLor7d71tzdr6ASrW1Bi68lyeZ3xEBSxpCc5BjI
v5G+isWECFa31zgyZDk3kI1xQy17d4Dr4MxfPeC+AWJp2E9HkqEHghUEkYap8lVC+KUm81cFVlZW
ImJu9wmYg/QbQ1DspdL/lYCyBGFFn8xGr9vDw40INsA/1CFDmxZnitRRp0+9Q6Vqe0ESJVnHw85y
mqUbavuXsUtnudhhJeFhfn5FxK1aNFnEMGPGyu5cXZAMRyg+JmRB3FuQHBEKh/floGu2Y1705Kfg
QRfUUTXovxwarP9NsCBuH9pNtP8ga/HpQFIWg6wYzH7xMgVqqbbcYOPF6u1cYupUXP+8UXGYczuH
mVD89v7anSMNMCTccvBq2TgZtWzruyeF5LC/yxpp4lNy9hxM9twVx6N9fBh5SasJxCVuNyVxPCRf
sJF3vi+j/VLHk+Ee8g/3OyEs5Lyauq0XsonpIKXWA6lu0Jj79uYtIItig0rJfEBcZdk5VQX+EMZ4
vSEUrTFTs0NfZD/vtPoKzlp290J4QpMMRvjYC3vmIJB2Jq4/i1JjUgS9+dSNjjOHIE3UrjCrhxeR
sTBFSTjrEgnkJcFVpN02juY+GMThcNBGrLv0wHn86Gc7tX5pbHv/LIZwKMFq31x5Y5nlNQ+pkfgK
jNWIn+q4Me7PuwDQrF7ENgfRIH2/jf3oEwX6QScy4qmuKSvgnle0PFMRMokPLdboYwyoCit70S54
zYQRcXxFSt4xp6hvb70j0esqeiO6y3HsHwH6xXUuRIomRvfrnTuDbnItF39c8SMFklxNwWYBg6ew
30ytsSB6pW1djAySEMS4SpXrVmtwMSiN7pONmFPmd12riXSvxKFgOedqpfg1OvZUjv+VXoldIxmG
Gd9diptMtk0PawZkN8w2ZFPnqKVa5PPypJVPTttiGB7qohO/qekIkAhF3Lxelj3wpnoMueT+Px7E
Hi9MpGYWcMuZZxEOGMN8AnGfdZpIDUKTU/ELBtk1KNvfYMZBFxZQVNT6HzDg0lHWFNnIhyXoUvwD
F8aw9Nl8lV0Doil7eeILhBMjKojbI3QSjsWXGmdFZDKyZ0SiDH4fAa7Vvy2XLtaQLGrtmV0yZt9H
yeiAdb4JKcX9K/NAAXrbqlijYBz+zqRJHUmrRTDnblG/GQGTOlfV34SnnHcSu0CMziWs3CRmY/BN
Lf7bXY7ZG0VEBIvvH1D28x8aasAWKEhLwb9klR9BHTY8uYmqYnrPfSRHW8qYtgyaNJPgiZfB9dDJ
iuElnwb7MeaYr7wP3PVXdlyVNgydxHw5gd/5WnzNL53BTWC/D74rXY6oZElcPsRzfFjZY+89xSgi
ahxzLfjJaOgFHjHvUqkGFF9xe0jYQ8ujPbUGdxQTeYYtUiZkqYE6IBY08cgldXRMxZCrzD3FfIGw
r5md9ZhvufKx8V70lrkMUEHHam73zx2D/PDrrM+rpVMZT1ugHWF3YOnf/pXxocSxUWXCHtMjT4ID
kW8mHgxFFUlEn0NIKK2yYDky2nPFGFfDS3YmmlOjtRakTw98kCZlOIpUWtb8A+VfwimgbFRl4ZN6
ittVR498c35H6FFSa95oYtLuO/RTynWsbk2p0dcutM+Qauil6U4wvvygXXaftxra6bI4K1b20iPI
2X40ygIRq7yPDNw+AAYYAXa3BhI/WPw3KHylsVQIR3nyWsm8EBRg4aGlUBQ2XH0cfEeeuk0sdcP1
MRqLSwL/L8zmB5RgUYKSkCI2wA+Smr/mu3ebp+cMZrUrHYlsfnf1klNGmEuLQ/dTjLFZoCbK5rFd
SJP6RDs71Xq4G3qg/1/1Ta1xrJ8m2u9QbdWbcpsXUqcaUi9x/4hSW1AmjUcktns5PtQfUnGO39Wx
dFBnZ66Fqro65QtYMdKKkuJox4Bu1ciZAK8rrlNJ6I9Wt/0mQsIXPFblYLemB9rOTKeuobaxMhEL
ksL5YeoDat1N2Ac3WNFWHu71eqlBydE5rRkQ639o/YQ+Q70u1ZtyD3S+LZb2Do8IhhfkppS1eVN9
S5t17tx6/p/f9w3vyxAyOIXXlvSanJ0hZXHrQPrEZe8I68U4rMRBPwTgG2uNZrNC8rFjOdSWU4ki
gjn+R06+MeaXg9xrOCQxcKBw5304ooaINm4m0OqhUrf7h0AC9gFj1CKBrS345Kz/7BsxctVp9pSA
XqbgtGHenMuSXlZ8StjPgR2QaUOO4f5n0TjlIImaO+AKNjkhY5dVlrac9VS9HHNtfSxkJnNeu/Rv
OYLN90e0ZyLdXFUpejIQDspX15iXj60XnZmQtNzEGWgo0N6bJcYKx/S23pKqV9aksQZBBVvpFEnn
wVtbn08i/7JvEeH1Hv9f9YQL7i158gNNqy+Vzkr/NKF27sfpeDE1+5u23CGl4S3huZF2EVUSRXN8
cy9bfBRP/zYx1zJQjow8eDsDotHAlexNI4ZAjqtmV/zbxQmAgqYPqFOVnaXMIa7PK7JxUat17woc
Y354rd5es1ttd1JX2UdOGkQrew8b9yUmG5amquQyZk4O4KrymTM3uucWarHDJfgZ3egnv+l4fwjt
AU8GRzS8bvsUQHqswsq9Sl+2zzyvYxo854VN6KTzCM6cfhfiniO5oJnLrdEaE8Pvgy+VZMkQJayp
3pz5TYq0q1OO+RMQgoP/sJxIrWvnm/MiQ/r3MUTrduvosc7iCXXxEbMTU1I+ayPC0lAPEejeGrd0
d87TLYsnOvM1XEi+kR3YIuPCPzu0TCsxyjp/04bnr8seUAtjLXPCoD0jvKLetTDlHmoFBVFqlCXp
+tP0kNev+XhkHnFYGX+xFMid3tMEG3HxXmfQZ1IuqfOFTJ2JrhZHwsYaP3zMbXuXzHvfj1qfsjTp
/iLsPnrRxXzUwVFj2wN567W1OR2xr16qjmrF0VZe0QEsFpLo4de4JT8Z2yTkW8PVkNKLLfMBunyx
pIAW/80H6Q6aZtTa3IACkOZvLvQhaFIPoOodgHi8EwJDWUFoTLav+mpKmE94sJ8/RkrVrjEVXrhs
7xVo30tUnM+7pKZK7bJLCaPooWfIkfdEGPkwMX6wtgL5rIVTO7B8eFdcTYfUHP+sSXp5tWMr8Ieu
Hu1/zjvB42uM9yu+/8RKF1WL3w3kMpgMIMG/1lUW5EkM8rvALHNZhPwusaf6L665V4SwZ2CjxTtS
pVQIVnzUupxgsQ8/+uOvx6BMRUGeJgr2ZzAdeTxy2DzSxUXfhgqLYMbfkCuvMApWRwmrK/DK62zo
Qz77L/ztNShZNKPzcU9Y4fE4JHXpv54LMIQw8DtJliQ9ZBTPIdOomxckb1fxS+VRNWjNIMYroj3B
AcMNG27SoSO72DfN+ZiCQ22CdG4Gt5tjHyFQT+bMaSc5HqSNOjxOj0NhaEZbcfDL9TOMHjPBLXj8
X5FPwqPwX+JTEh5suEero5z8U8v9FYjy+3jG6Ly/5RLfis1ujrYBTpIQASuy94h8toghfiovtDL/
giwCmsA0+6B+P7ZE7RN+YACAfZjeRJJUMeVTBx8Wb7RmiubfS9XkRw70smvNrIwQ53VrVbhnk1bQ
Vls0QRBuQSVKKU+gPJkm7PJpIzB+dGoILzMONDAMIASY8ARYpBLCRPJ4q+vLtXDM031kqLWWGmhN
jwE4+RF1cms88oXwF0OIzdv2A0phQAV8dOZ+4mDL1w8J5KX/whY7zw6ZqU+ZvIbeu5s9/3MaA5sr
bSOmpTMiIKreEPmLS1gNcjc88I10atkgkAhSnBn7GKKg3nS9ufyl5QbI7ZJ5/HZ5ErJX+HUc5ADp
teBZUJ6Qdp1K+wyEn2YFZySEuGZMCwI1c8E8vjm9ia5c2LbHWqffZW2iwD/LPV+rijlPFKHqst56
fpeicA+Gu04E1oIf8pETYn0+zJYyjTX7LSYK1vMCqWnvC+G0zedNyNwT/DDM0DtgJnwEeUp6AzFe
sw0GfcIVzanLgIUHvk3SdNEeTxh7xJiXp/Mb5XlvmKz006TVgzfrV5iLjiJGZ7yxRmKA+MpsIOvT
TeyJGsCw7DvsNe+jfF4NwzbcUVVAtuAXi7HDhkU2eBKBtdEm17oseIAFiYd0JURX9wvKn/QUQYJi
Q6xyZHvmxSgvX63lUCYt5Z6rhnLC7smiw9GXqjaAQXauLBkIIVHerKnq51bay9MOF9lFE/ulmcYN
Fv+/FhhMoCnXS4uwcI6rN/r0EDw8fw/xe6KTWRsC0drASh2gc6aCEFi9S9qOH6smIKgIzSY8Nq4W
xublZRRYm2LSAwEeOOgEijYxBCD22cLWk4d2so9umzWKQ7JodN+yLVl6OCifn1bHJ6zdDt0Vgn3w
QcP0C6zZgELMd9BAM/qvJD2oeEnWM8vGmEKd5QcZEyrE9me9mAEKs2g8YXkYNHmYJTfMzJjskdgD
S5ONlAVWkNd5mzkfiUhrJxAGRIZ4FIQv1Npcn0f/Yw3fx0PlQyV2mu6/24vILH0l/yFt/42YxHSD
6nMSBJ7PamsWRrFcZgyp27R+DWELNziUj6Q3oOKRctD8p1wT3TSJL87Sy7c3c4m9KROx0RQhulGK
Jry7C6LcGL72iwqcJq6QyOiLGSwOjSJckn9bTQVkLxWurvTBZ5xDDNNVkZBwnGtenlWvMJFckxvF
mwppr0jvY1DYW+M+8iH/IkrLFFnNjGdUFjrQL2Rfp7Oslxt8j81A/QkwlkpIoHODGRgB1rSiHc3j
0xV0VmkfhihRrYuOu5s+wr2D0Dzi2Id2vRvSR5c2396Lp1z8cTJ6otOFz1e0JA5ZNFz287uTETMc
0K8pMXtjuVR4gJ6ZysY+96wrdB2vkUzCapxo0rI4uyerM4GTalCrv8xfZJLJaebsZp4aJE3JbITQ
ZEcW1h8TbEp4Z5t+F9ep+Db0cI6I2YAqOKp517TNdOEQJ6cArBIPRVDJoV+1lGKexDow2OeMMi+y
EIJ849V9G+Feo94w4M/Z+yEBGNaOUf8dLBCeGrk4cw+DUAxozngP/b6Do/Jdjyg8cyB6jXC+0QKG
hj9SRVKayfVAVFru848OEv6JPreoSRcAyBYOSPR5KldFGKAqsjUy2HckoztPYAsdeIdbdt/ve3Q/
XuIMDoNarBqF/ObsIGeWfNF1MBvun4a1CqNXthdNf5k+9nz8bL6F5hOHGsJC0RiE/EB8Cx5d19S1
V/IzCw33xKLAjJ0ICF+RyVYNBP4xWk2ZPpah3GI6jg+lSacnHIXAuUHvjJlDnXEuETkPDMGPz4XT
PDprIf/xs/n3+3AUruA8eQxX9Yoq+ZwWHLUtSyCglg2DDx4IuHKoyki0OmF8s6GckpJ9iX5nG4aR
P3gFtTjWzxAbkthVjtlQi/WjEssGCXD2ey32R3Dril8XaIRtSOWhS1nAEIANng0x3+m7GfxoqKeS
GVEsREOXfjKeg8UmAd8F8pmcEydbnw73/dcxNjyl0b0Fov7oXzSiqFygMCpBM8tI12trW856Wipx
HrnfAJgOZux4Aau7VDvaZh8Ml4lIZ/e81Jwh4h++GQfvgaj3OmXTMo/I9XErWL9gIEZyty+DvUiG
iCZXNJJ2Y5WjC+4bZH2lBTT4Hh8G5NWEYkt3PlPT1xsCr13HE4DiY3Gy6CeILp0ys4FtBbgoOaS/
talSZIDiYde+tRtTuqQM/0TekPVb7Cb4Pl/cUyO0gZqVj3sLucVtEtojnD8lM3A9j/4IpfNDVLll
/gUEUIxkIsD810PQXgM6KbqbePGRKEE3MMU94GRCx+4MgFgd5XK1mqD6EPmT54Yf9a2BTf1yF7lm
tyzx6OaZTWfCk93LobLGJVBli4N5A9TIstQyH+vSZ2QiLo1T30cL52OFQQoqgohWAiBu+fFkSgYe
yStnUNn1KaiLVtZzi4VslZ1MoIXfzSlnOP0lVnuItJ1QgRuqDMoT6UdNw/QC1WUhlGZudXDHvoqv
plKfW1RGlGGUsQ7V5sR4vRXYcK2uERDcnnXKbmC+4a9mm8qivjSene0nXNogZDuLqU3eqvPNIjO3
cpzrtAo5vUeR3H8Df/FXOwgkSo7xmds6rvTYW0Qocs7INAtPcFYpvg/mE9jftKxMOJy7STaoSFVf
eOmqgWx7Vw3/mgl59mHZ0CwBHj2lDAuucEXq6FEY+Dp31c2ltZeuRBH+zPcsl2DbwFH7/1f/ePVy
pVr6JyKKVyXr8eSIUn52BV7+zkH6j48rnjTWplZtSB/xXNFgol0Kzm4kOmAg10yrlkX2VzCNp7av
k+Tvmz9YvKGx/jqIyfN8sIbuHhT+yysR5ZO+RKIWWVlAHO6geM7geij1WaVUf/UPAgn9ifokGkBu
n4OKc+c7Dc+yylXtgjFftH57j48k+2MdQK1TIs+CYhcn9iOhN0DnmTZ7eBvGr2UfB70c+/6uTBV2
sGiEQ61GDft7gKblySzvtFDUGd5MQwLAoPPHdef+6Qi7SeEMLt6BQhMd7Ekbgg1/TqqI4VIro5NI
EGrA0qscvBmnYvgoXaXVenLUtzfd/6OIzusoYKWzLH6gb9cEtCNJIcLlAi+0Fhtt5kQ6wDbZM/Mr
CZ4lYsa2SCEft79eG4kdWXO5CHrTCvhYnMF7fetG70vDh9zQH67QakzUNgEfvGaF1El8D1iBfoL3
8p1U5QmU8mx14vcGS4nKAILvR6vED5jhZcyvqXQWukak1GFHNAYtSkSpt6tNHP095epNUOffpm0r
J3JFeWS7yIqJs/nexSFy8ER7qW/yNkcX5YYv1QfWi3k53aUvUTi7tqqKbVrXXD4BUgxw6p6AVorZ
YZXzrZ/4NRaACq++MmTuJZs0J4ViEHWvrSg+C8NMEeSs/XSi74AzaODCnwxesom5emGZYgKa6z9i
9evecSbjMowLD/EsQOfr9gIUI4wbdW6hK2+EU2vzHgRhYgA6RbxdOa+6FK1Wsp6gRGSsXtq/s60N
tm9ICLu3uAqEq9KgqxOhxosZCt6DUdBoi8d9VC/eQq0cjtiY9YDOnuZnha0Jl3DvbIzk4KG6IkmQ
/Dvzhw6g5CuF2qHA/GVf5NyHRguK7XU1cnYd62qteIS88cGArThywiG+vswpiFZG2dUeSaNTPmNx
en2m8OFNGY5SytA6tNKECZBDV5/xD3/HmabjNw0DPiZaIthR1AGi0luq1k4TX0T4BbS4r2YrU9/G
x6G2JZcF8+gVzMIVmJkpq5ykwdy0vXCG9PQsnBR6fDJbwQ2fsWxPxnH33+2U0INpZXdtCD0N9NOS
DCXpdOhNc7QvkL0c1NzfVdEIlFQHErfNdeXgGeVKyUA3DTzI8VOTiGemzgFQ9IFLEZWrmVb6ZDHm
X7r6G8E6xXK5gPIGqL7Eu9QUfeu0c5S+lljXWtuNA85DkfuHBLIKbCabOZZsGERBxuLbDIzfSqHF
Aoh9kSmgt88FyK8rc3oWUWDAxJDHm1D1eniGCZd83zHA+eQoUnLLn06OrcnBlj7nW6m11LgQYcMp
4eeFk5x2UJfK4+rzfc69kUj9CGB438Wv/QyBGxkW7lPcRaHTGUwC0JnxhOn7XJnBfChAC6a8FyoC
jsfc9nGqXqUIGnAHAaI5XF9qUVDT0w940nuOpRa4mPvwWIrQ/amJ2Tb0Wh41A+pQbiXBRaL7fwRX
3LEaVEfDSWziZN7o+gI6N+Q0VYxfiJF086Ust+l7j4jPOj4vzqRTJGf8t3REjUQfUUCBaOtPAfWx
d8sLR59JmqRI4ALYnfeh7Tu/GVig0kGyyd+IGq8M6UPM0P7DaCcM22gee5Zk86IqikPLYhW4foy4
kR4+Z5OzxDn8Qyg8Rf8LhLAy6aRPwFpZsrrrCb+dMEGgheY0a3iBYcQOAb8EFaSoDuxJE9rAEziX
9ncWO2AKkpX22lQX8/vaSEUYb73eI53NCKGn94hNo7qqjhBfuEmqDb5x8mT1IUUpN1U0R90nkB4a
Dyna2tC02Of/+f7JfoQmjq9pzEpRK5IcLGdhMODZporVLLH/Hmm+UaN4Fuajw88r4OJAZcsFHImb
CFJOgEwuVMX/3ErkkFg4mvhNOSqozv8vdBttzfa3YHWMGoMDa4hEXBkUNEI2cyez9i+xi0rp1Iya
FO9e5GmqfeVZ3G/7qvJdrF066+kAR4cFxhuT5WV1Fa0JSJVc6ffQ1jznnGNyXkkj+7Wv3a/YLccj
t07pPCRNIeveEmICvAjXDWsoy/NyYxkcJSOtLzWgClVfQ7w8M2ON7qhTvOxAvjWt0Rv26R7sHlYM
X16IYh+RRJOPurCUJs3XXnO0YdH9Nsk7Zo+Jc4Ej//wFqynZ+oNIk0JX+5loA/Ht8Yh6zvLECxkm
obuenP34l34J+9Rm4E1n9PMu3aIfu+DxCa1yj24OHy7GQ0JKYEfGbC5683ZX7lXfLfWgQpvbs2fo
0fmZ1TCoFCNghBywl+JcdR8U8OxCemwbAOGMIuCFlYEOdJvz9K9Yz2gcLca8BaSelfAxy876oZZ6
Mpb5TzzjdU6Rd0rn3y4oCetS7bH9p5RgqKjbvMA4utC94lYACFenQicX9f2vM+z/2aEQwwvEdcse
B1opjWB2Ax58HUy80X47g0ChF5pgT8jkD2f4Fse/1P1yIoSOk+d4FYPcfy1j1zokGjknYu66SJA2
xs7x/Ns8gM0PX5QXcwgsQsd7ukvv/LdqAv2vemHb5TiRNNIgpkxbGkDqZw/yn5HaQaHehKo1M/uD
ei9xgHlkjeSchgAI+7alLmdyfSDo3Z0yh6jqYqJzhPti1NSYNaSYAThjUaLcV5DyzhOt5Y5683n7
hgjbCxUh1345ESPwRSH25MycciDeMi+YdaT1r63I4liRE+DBerJeT/3/bCk/Bq+/d54NsSzVQj5b
6yaw7HIh9E0CGT06b9sRYNc8XT0jeeP2jtXVNVjXg0DzJBJddumyblYbPzQL+eIwSJZA8Xbdec6F
ELpITVi+y3gNHgUjMPK0/ZYRKu4f9hwXN61c2Jn0LxGzIew92o7XrtQVGHYg2nT52CUPAa/bSNDb
VfyBxPrhll5iiJqG/LfpUnZCL29N3ZVgcFWCRSOBOk0H8eS8qMzHao4E63l1g9t2vGx/x71H0Wzl
RFxbC+knG1j9OG3ORljCZKcCF2mijArADbHJ8i14tuVR6u0GVhe9yhy2ExdYSwniyjl1F5S5lLtk
qREmdXqMKyKirvp4rTCeOPWzA93igymMBLivwWYppZpMynLCit93CYBrWhBdgqY0ijEAcGtYYC5e
HWfDv1Q9EXDq2qlt2pWaH+cnS/SdS9tEZy/zDBAP70eCQs3rW7lfA6ionRjy+yk8gd70kU+mrFo7
70tJfoDYLymRC5wHB9Pd2MBuQuOH2GCoarC0lDQ6E5mSg5C+Ps1TZNPnM8c/kFKPcUwSiZv9w9fN
upZwP/Kq+lG7dGt+M4EgbXeQg50MAxjIOJdTZ/TerIKjqMQlgAhvt39PMRK883b6cApUuTWLu2lg
72yB0mEvdOJ3tgItUPRAD+XY7xyYFcfKaGDMtJJshOThiHNeZ6bj7RHerQQM3IcRKN15AhO+xUul
RdqJDo8teK41/C5wyatjpV6aUzvqjJbJA3qvj851nM3N2QWpH5AlaK0NcUORFjMxkc0S6vtkTSpE
+eQ8/ges6UDctqciX9TlUUZ4pgDhEOb0XYG2Xqlk11opurIXPUDB1Sh53pjN/x2NaOju/6+bTyxv
g2+69nygyW3yoyTRu7noYZfmiGdnCzkRa8lM1PJr6d18iHZ18kICdSE4aMeTWWiEaqM6+7AzG0AA
eJcrjWd/Qa9yZUIix3enaZYtGv5NtMPtpjHR0AXyv1cs0fRcf0Sj9ZXowC5g0ODHRof6n/f3drNQ
5w1SKXZDC8K+CkTPKBSsO1R4cY5CPDr7vrh+xmGWq5sqDUa8ZrcCPxsX4Ay6AgA/35W0kgaX3R6/
kZiPd3kmD/6Jll7UwffYYSSgS5XXlVctotufR2rfaRC4klJhp4yO5kGdubVUBLNPzz+38XQPoqZt
UXqeiLnl+uoivKZIJZ1rnkA+LxxqqGkMATdoF0RkA9jMcSCoYOS7dUNVCV6NnD6NOza1f0FlJgo2
NrjX/JpFuj+EQzPeQmQuG+BHkkDxr0la7A0mcqdOW/6MGeS/0s38bf64KuEoaspMEJD/dvG66ot/
FilrLIyZaF7xmkQGS8RKGAv+KeJlLvLncScYDdLNFPmClkK4gW0Ma2ICxyEv8OkfAqTstitg7p9K
ETbfMSIyeF6iVCd0bqR+AROdynq6bbmGPGd5htBXoXE2JN1vJefSGtaMgXlRfngCt9EWRx+Xx3Kb
AhyhPiu9dtPrJGpVdJyzuQvjdPybsJ5Uw0s+rlhDQEKZiXxV6hl/bKMf7rwQf+5xUvjpHOWeq7hS
ZhJmQZiNnNGgJujsV3CynzoD6UGNEQOgPVaQpWlaHplUbQgfKkaFhV9DWL8bs18lJGJO85BU88k3
Qk0+VKY4IoKLJ0A7TMLKt0AjOv6YZooG3LacBgdYfo8b9HkN5MJqlwbafzF5pm5CchG/G+V7fq75
PXp8IYkho1i7aQvLlS5ufjdb5xGoUB1fUCp58WoTu9xVpRI+Bd0Z3kbHckCwEmwejTX0cP52WqtK
DWPuM2ZFYvaFd5k6pk5AqZxYkILMS5rbze+jjV7PTa/4Bu/DtEvUpSf3CI21IDl/n67ioxGBvrLp
hFjs5H3CANFR1YVbDD60kdgQiuhwPmo0Znb3I+KUsRL7djjfiP5QW47aiUixuB+hlm7bPuWo66hR
O2OqrCMVHikNdNu/E7RCZpuCSJwCpDHCZHUkU54JuVSjf/f9UrP3+QqLQW5obQqXDJCRZ7HXOlMA
z2qjbmIULS/nbx8cmXh7rhOZ6VYEuuLjzuqsjpIFjjxXP0pRWvoI+ryMBO/+Pt92kB4BlKSLxHun
SUuBaU8WAusXwrZDrQracKxo27sU2Hjyx80TOvZrzO5nz134C5w6QUYpMCi+kyCJFDJzXw+osGlx
qDk4fN2Xr1aafCoCNkDUX+fE+OiH/fDQbTuFqJPOjmjrfc/uoulGEsdq0x+7rjiAuQMjIovrXX0v
H3/niKT8IKUm6C8idg9mcVzrQtDuyulgFYtQpM4FhUNOz/nzE2BvJlYURN5exPAQpjXdJGnBJzfN
sKg0dVPJMMlcg3SP2iIYvgSz9olgYV5fbhLgWNnYf+UWO1PmXEX8KjPvyJ9sjcAnkHlwj1qmBNPb
t+Lx6/4bb90q2WnciM4b1fMLt5Fs4nuto9OciSzxvZnxVRZPPU4EQjUzS4jwY2zPln/SCMk2y7a4
xh9xH4q0m0IMz7wPAIno3PPF7pyuJ/4dYN0mtKFQtp2vCKuPx489zPaRZonak3UaZaILCdPLKNJi
0M8jEG8eTbmdW2tG+rzU4+X1BfrnhbbD+3jgRRTeUlatMTB0av4Gvqt1/wUUI55PKhQImRT24nI4
jRglGv7ggmw2rsrUWoXejYSaFsB/DyvnmNorT5k0WtH1zM00LQSz+gmaU2CCkhReHUB6AJOEdhVG
SAfmMlQWE0EbnZwdt5fIGa+LB1yU8Sj40V1yLu/qChjrCl1HPP8HyKMuBLBuFRihUlJrFmlv8FKh
37Y0Penzy8RlG5/2Cyl09jl2fmhQVG9rkEd9dHVglOoQR744yc0Je1o32IiGDOUuAnRZyyAOoFTq
mv/aKAJOJzgPDJnDmp5ptPgfOe6/5yYpgst0mj3h/i4ij9QtrlyWm0BnKkO6Y/cFAPtKLK26IMFd
qoc4RgejAo8lnvt0DH92S3aCksUcDSpZIdzntrdv8bPgO4/PmYeqqKSvfruNUCdKBj/C1Vb+eSr5
7gpMUkvkQrtqYZwcNjwI58y9czu5EpCoiqaocqWoMJJcEbx+jqBp6vFdvtHNHmwgE1Gbi3wlGVfP
Gr/tvH0JS9lrf/J31shGu5la1pZSCTyO3sJRBCrrPPJD4nr42kzKrwYEv8SwUsJnDBg84UZ7EKEJ
nfx6Mqd6ATxfNfEeFSBtZuJf5VQ94Rh3Jx98RZtsfqHyjgXy4mLKuUlhegL4Gu6oQyPeEqI3S8db
yyXJTRvSCDSjqFgotd6g3GiHitCWXlv46fsXK07jp+xmkDBbsupjMvLfLT/qf4LLQpkQG4a/wVcO
YzqY79r28TAMucQ/YvCcZYFnpquisNPZHYNFrMSfdFpPxfmOiuaeVLisbiN8R1tbXnUDd1DQu6Ei
iRhdmbpsBA6ZmtNWLkLg2EX9WPMXHMLOVaZVp0fJSOms8bCE0D8k2oKmTB4n3ucc4j1uuNf9J+g1
KFaR0cN52vvmj6ueheKfxF4xeN6N9nRneJPang+uTLEGcyMFtUl0R6u2CXoQ8OaJePGSRJPeUof/
iVNloSafXIkL2mZP7RTq1DOO8BWhl10W2O3mTyJM2D6+l0VCG7nquZYNpAOm/RqU8waldnGzDn4L
FX/fP2wrkacUUUmKpDodVSgBTPJBxbNDNC5E380BLvBXV2y/TkgjVQh5hdUuebg7xqEwmHxUjL3j
Dy3o0ZXwJ2lIngovs03j3LU3eEnp1+uvUaUu4EFxLvD+KLo1JZvKDlpu8QKBNrei+p7+DGG/uLKn
ZvLQ5QS8B8CEQTeJ2ehQtYsXgGzV8YekaR0ov2eDZ7v6QOawFcYDQaduaOATUvBXyh+jhfjXGOTd
+vTW4sDEWjkv9U1lBx5a7q4k1ib07VD+8xmi7EVZFejjaXbVkesDfReY6YqNcRZXo+dlsnhVAE3J
rf045DU1h16ojvVXy0rriidKB6Csr+Nhk2Wvi1maz8D6c8Bw/HpCAZ15xYzcXpJE8sExmdjawcy2
KoH4WhllodiTbNrNezsXiOs9UainLgT3NBd5KPknWHTbntjsMYVjRHBQ3ycEHZb8y9aUAQcfqx9r
JMIExMQ6ItDCmgSXtdvyud48drZbwrfCNnKMiWbHl0X/yfHWcReChTeiIlfmRjbWxpuohOBZIx+L
A6ukuoU++CjOEt2OlMwpBXAtj8O9c/TkJw5qSl0XkaGNeKdcFSYhKwy81AUBCmf92whqmDWfrjz+
KDayKuXM5/UlIUAUQ2PlLqmZbIXdseJldJr9wBsKDsp8WtWVu+t5pJ3qnHunM+7QzMTu0w7lkmZN
b5I8SF99QaU8FbEBP5a7PUevc2nkZVup7KR6smx186O2x22P/xLEtNpkUFB28vLmsFkJP4yY01lm
2YTiGpPjLQayougwCEYMldbC7uZUImcRLFVK7cP4g0CrtE50MjexDqlfQlq8EK98nQ1sefSRQW8u
YuTX1oxcQu4GPUqqWGJ0YbGihUCdxZV19H6y2QZRdTwQdba/0RWvNLKDEMyGCwjZnZDClAFMQHZW
q0FMw3Ck9RlnRt0ZU1Qo1bKUMnMH+uZju8wNxeT5uviMEawT3qyC7vw+llGLGiREHidzARv2azQz
LE1vCnuJD5pylQpttflX0oIE9XcCRfdWY79x+Dmfa9O4UWmwh2fRsAc3dN1e4CQqVMqOVzZyNotx
uE/X5nzwE/4vuGM1yMywW/xFrwyN/plzpbf1tOQwnxyx50Cywt9S2s/F2bYTQuzn46G9CEwoAoWQ
uafefZJkhTsBrdB9a2iiFioBBIlHI89WHqq4TJAOChdoSXbrUzVGuZBsY+pTWf0AAUsPyxePE12P
nhwBAXs5eZoTwkRDxMRsDGgwRwANRYMgkTFm/cevzpw7MqzNAQUkpMBS7VJTMe2LCv4OVJWyClvQ
Kp0Oz6Fx2w0Mtz/CH+KgnP2sWdh7fFrz7Yj8NVkWeKf6k2PWAkSfkIX7mzBYwaMwhR6OhW0o8k9i
1FfesyxTPkEctZLiu4JxIUGx8Hcl+38J8GLZm5ftG7O/1/ZSjMOUBWm/LRs0kUd1GZVFvVfUzLua
WiS0ytHa3Ehiivz9Q3qOuSE+Eie8LkkPM8dOq/SJS3OUvVUGTPmeQgh1iTbkXusHzpUGgcWMRz4W
60fKJYpusp8WLGUhMfznMF0tHhojnHv7VBV4LVfdF0ZQykdvJddawJtM+a9cSnssKm21HNE3F5gT
1hnqvYcgjLyDJ3DptV0nBm+vXN4Z9GHgz37zbB5eU8r+giKqJFBIXFUaQoqNRdwTWP+gOBogcrxS
bD97fVy3hI9AW7L3X6zMvmXxBsX6XgnAbWIZnWeLhoeV4fe22MGlOZABxg0byPTtXcRZ96TJGTrE
AZ9zFO4zXDN4yxjLBI8MSjttZBGXusUxQdNE/j7Uxx/0NvG/7p08Rz4d/XJlQ2983dWCYPWC9F+L
L6e6OSL/scmU7yvmg6gh8NbsRnpH4HuAIkFPI/sp9dSC97u10ry45utFKeWLVhBApIC0Ps94Lrsf
8/cd2mSypS7JTgGfOeEeD6U9hz+hCT9Ksw+LxLUvTR2bgOF2CzS2VdIc5wuaZo3EMmYjA0r3wbS1
6lbCeCMUdGWCgEFcJjTUb86ciDTkeWJOexdTRZzKa6ClxonO3kO/YzNcar/TDKyWtS0eNHQfxG32
4MbRxuDbGsvZ0+gLZhI7tq88t0Za/rYBxz5Lgy8JxLrposcvhSJLmBndQqPRb1RclsmN2+mMWkwA
HFzyKFry/sgAe65oMRQ/YBhD2tNLD+xJmWcF835RnkMT0n6UlXbpdrJqWKWXgh1qEBMFmIM8L01j
I2X9edIudoLw5Mbk/b2SvuOUV3aBcrp1kXWpD7lX0CH/WXjzVhctnW+wOZj80OcCchBJKgXptB+0
PK4kQKcCXI1cs9qKj+75wwzc4/6RVNjJ9UNCvkBMN5IjSO36Bt6vXVcxf+SVBKCSl8NvN9mA2PUK
kQIAaartX8YhHw9mU+au17qMy9tEHc+mqdiSv9Ynf4ORW8RX+Wjm8SvhK0EsR76v25OyZV3MUJmj
Q+6zvi/EBxBEjqHL5VA/14fKHCQX7HTJ4KuKJ6u3NigIZPffONereMwIJIF+8akl4K8br6AdHrX0
j5TqZHUEdzhnHeC9mS1Zi9c9amsaslBWdg+umf99ZmoPvglxeS134uHF8a0jx7WmzzHOfs1VKJSa
2zqzaUteL5ICQrl9jIZGp0vG3la6wQ+8/dsn4b402cmpmutfFfgSk2/10AoDZBJEvDbtgoqAM0Kf
tgzX4CBRJYnc18DtWVNxJx1HB0pabDhjoH+TjknOIp5i2P3o6FLMhmQ0eSt+rIwyMXGt3QCnNvxh
l+MfRQTh65d20Rls1oc76HyZ91JgNwUbjj0/gNkNl5pSrKDtsJf0XUHIBEO0kXOUoNxRsGAwzsRd
ZU76DRD47IVyHxFYFMuOPWpPib9rmibmmb3FifLbjMfPZHJ1GH5Y5pIiCsC8LZT10ETnzBPIHPyf
K1EYO07bd3/GjNW3qd+3DMJe8eXCkfnVMzYLi4Xy9SZ1mhZqcT6iImTUdrBWzH/1BUAeBFx3IzB8
wGnI3ywqtcJhwriivv/2p3HCISMhco2xfCZNFsLOFcn5s0NgWKpOnOz/j6S2NAQXSpp0BnJnGRxY
R1XuAEDG6WG+tEJz94ik5YFNmRPmjFnLx0DnjGnxYDEne1yh04Fg92+yWaCytx0Eh0MJRIXtcVFY
08WoPKBsFUMBWPuDzZ1ovmqWe/mE750FSp3ZBr/dKtduzFxSiihy1gwMIZuWlsfOdQMyCTFIDjis
AtovEo4wRKjoBi/9yAaKR9DDpK4ePBuY+wT/M6D2k4hTqgusV2ZSfHRr7pj4fZndzCDHeEdZkxGt
OeXtnjbqG4SsJjLbSgX/2Fbxdy71exPTuQQVnMGcgk9ffT0GlUgKfhmGHx4z/v+HF/1M81ZGRkoD
V2w/qTVQBprjfhP5HN1mTf3MeJjT51cwtr+E/O2hIMbHavsmNY8z/VaGMu7SqzsShRoL8aU1dgg4
3qTZprf/ANQBWIZurX2mNDwmkqJr1tNzNTjOAgzxvaVlnHIJET/W/rM2YeqGTg4qYJZxIyPb7Jbo
G8wEMdbSF5GUoOQcaEMId5rq+EP8XgDpF4exONDebcxikZQVlBfJkLrI7PorjqpSrzdgwaVS0Tl1
mk8Af3uUVFJUE0b2fB2XB7doQ6VGUC2AdstYLhiB4soEwwdmSfTtqO7wDd+VmXmiBqjPkCr/txFj
6hQDomfNRz/R8kwJEtoLn7lPOS0NBjXCpwJXNRIXaE5bsV1Y1GmsV1z3TLwSkh5ypWhkoxeo38NP
GknvcNMokgcMkHtBm0j/C4yW8EBK05CmFu7BpDnlbuo9e+crVcl/WQRISAANqBuyn/4XucQcTn3W
8rk8F6JqDa586nvOv2A9CDe8Scb+NHotOccNgRHZq4IcycnrQy8O1Z0vEkPhZ4p1hHHGzrVj4Kby
Y2jst3DU7vT9eBOLl7lxQ6PknvF35AAGgAAx0RRQrSKuWNT7iKtk0ID1p60SAC8CUkK4zsf8YPTg
8FoY1JeT2xrmVqMD7to8HsHyUe1blVU7Ga7FBtASQgFLU4AlKAnBLJYyLO4MmiM4D8FPgCDW7enZ
6l2+meCcoMTsOzwcf4X9EUpgm33IEO7uaobWnzvxjEayWelGfPrq4/+J2ZJrGw1qJ4BvbVGt1pu2
3R5ex5yhjDf7MUelc3+pqZiKe69gmbSTTrRw4ZpcgS+w25CnitxBZgg7gV8QrdBn/GcHcwHL2F42
ymwa0fTwBM9KcKQX5L5uQ7a/b2phfw7XPICdakMuHjOBW51pgQ6uAd1s7OlvmgPeSedyLrIHqAWA
DcDmxxsw1sWwX4392d6Y6pUjrWWQU5g/1cD8j7x+oxQPo2LJCBpB8orPHKkbbgnufr8mDHeERod8
3O9G7KcJRKQHflZlbh08X8DRm9PZnc2pD2zzLCpXkAYX3gmhjxy77aO7Hfbgkxb9EM/2K2//bnBK
c0JbLzGNrC4xZAQT/OJs33Jg+QQwYVEKYg5D2jvSVhU4Wa1F3eUi5Jzs8ERF5y/XAaaDXhrngKhG
O5418DtUxJSgQNGITdQBZ3aFR5QU+abuL8JsNYEmPUqSBErcy7Y9RljJ05zUFK21Vighr11lx1af
lSAPLJSsw9jgW5BSdKUTdTUyyqzA4W+/U7XIM7iEal3ZORcmJNjY+xy7dSYvOcDBEEWbu4NiXahY
XR5TQBMjmfSy1StH4x1FmJPP/liRj5PRIV052zXPh+2Jb2sAcrEH5miuLXHAfPaO855zdkBldeSb
1zGLyvuaDpNvXoVpkq7IkeWh8M8TU1wkFkqHoW+KZAIoPBliMRCEb3dvS4WKAzJzX62NT+8sVbXZ
q1uK1+PIUBL6XBg2IdtaFxX02ydNuUWLTY1CwqGAnQnVF/fC0JSk+YBxS8D9Fklv3/3Yn/1AFbz6
5LxY16tXb3CEaLXsXhhr936OURXiXhLS169FDRX46TRpI96e9/EMvznSHwdvM72jiYyXJLG7sopx
XupBVwV/P26xIXRtFuaXAeElA415Xa/pfSJ4IfVhIthgpt+Eq4N2uvO/OrLfmSSofn9qyStRW26/
qObr8Kecho+qM93vAp/1pG1Y/iiLkmyy3ztH5F8DTaMsB4nHXRKlSI6XEb7y/C7ISKN0HKL8IMJs
znQQPe3HSd9zZqFaswUmledP0mkJp3C/AzZ/iOYrJb/Tc4E/OdKTQXWOuEM2LhsIzMN1QEsSGVtM
TRpeQxrZIBiW5n11yVFSP00sTq58shxgy6YA7NKKRoMEWC3GLrhH5XUzNnzDW7rZi/l9Cqriydxe
7/Ul9K23vMW8OGNWlVs4aEcwl2SI1iTfHKvOrNNYGF6XCZC7rRtg4Ty70nit5KFZ/QPZwFsBEQTO
8CdEpo9fXJYJejTWXVO5PMX1lC0iZ7rB8bMhRXevf+7MQ1ezeRfFCPIy9NDgXP5VC81eT4VjSu9C
rmsLdfeABD6CqMt9sBtHysoU7ODkEnuIfGleSMCpEHmpO/lWOSVRWNCx8eSwAQ3wMULZSxk4syfx
cUhuQTTZ+QM3AWfM8PeDDFXFPHPfPwUm8s0JDUSz4zYxeNO9m8KJ/UZXgQ8qZYaOFJpDnK3vbNIu
tn+9Yk/iQXefMtzFjiHhlxa6mC57LjzN7yRSzJUOovKGkjUoEXP1h8bRf72iYmJg20xVT3FmEdWa
JHcGB+VLUmufvW2be9PUPv4TvJzWiGRjlzehkejU3NJtIjFYGakvk3+HK+wmeeCgwD/6/ywZNs1D
0W6Bn0OD36IZiZjncqpUdLA8d0GY5xu6rv0tW24Lg4ZVG4eEAs/Xxz9SW5L3gb0Hwt2UPz/0A/z1
2h3bHDRKx2fHt2VFoko18wryztGA6BGqXufyN1xhfjBu2w6i6tqWBpFcW5v5xQFZeeR6dcWEkTQ4
BYM9fOUvSF1bCz/FZlWpApqQV6is2in9FSjorl+EvVYUln1N3fXZYMtFsRlLdgnSbscu4P3UghXa
QoOmH4gzTWAz8tpKHItrz+k7XMMB2EZgjF9lolSvXVTGPJrgW5tLiQtKknLlOpDtg53JeJuFUxO5
Cu0OidLX62bFMbWLJChPZZlSUbxZbsvYqUP2BZBywHnzjIj7kKlScxU/wrdU+6lm+brjVcbm5fEz
vF1CpJXNUUdUjm+lKKYqyXwpD6wbsSXqVAaC2FavxDEdT3FONTcvjH/mBSgcbFHIl6JWMHxidZ1Q
Sm+1ZjfP7JUOV4ty0hbRr8rpfabNZ4pbqyByw+BxU0QbQcRY8V+btNgUOm46BfF7azBgtg1i5JDf
xbONyDtPktu1uFcppe5C8kfBcT3ospBwy7mBGgg0YH2DKtRbt+xmF7TupqwISGJ7yg7CU85esMp8
6yESHcvhDRqFxm0InStrn6AoSZQvh9Y9LMRYhL6FXIA/mERxamp3VFHmOvfc+40fpS2UBmq0XIUg
rkK0Bq+h9sAXBY9ssg/pf0OttF7YukZf2k1DQj4iKAsQwLq2QT7JGAbkjaO9fZv7wg6qGqJUq5yO
xN+WIwqOMvyXBARJfo9RFMWNpNlbIjJsA8e1FyAFLMJWMPZCZQhpf+fe9Ei9aTE0gSeW4rsCQjo8
UfqfENRnoBF6/63fCI5SX6sVBRbqQ6/iJsgBo/krpmOH0IPflPnpNc/Nr7//p5SZODI/W3NO5tQQ
pdJKt4t2V6bCTxr8prFdNpc399MZQMyAKEEMzeBR4RKWeFC7EWSBdiY/Lg2LOJtGo0GbjqHrWD3D
La/FRAR3Vn1odOqqGvxSIxoaRolDbtsgQdrJcfDfxldAlujhUy8v/t6qdTQe2fz+oK/HBBKXL9gC
3owxpFe2xY5h7HvSymjd2dRa8jTk7OFVunVDRxpIqRV2BS/JPaeDKO9WRmyxhxLQxF02O6X8smQT
llvFwp6nok/UefdWxODuZOcyzIQVReY1jg225cK1dPufV/XhKEfLeTwMYQA64vfyTmN4o0fo30/H
8ggTQtJ9y1gOAXOYEexFlz2cyXxRBjJx5dgVjGKphzwoTYqVTIwLn1rf3Wc67klZsjc2dGS6C9GE
jK8xdcSdMWxf7jhcZiB0GKCg5gAZt3ftQ+ufsyZp8wdVU37/yuZ3iVY/Mf/DmQkeI+suJ/R9aE5I
IAhVfbwFxqptDR7AJGc7OjvAS9/SnScvXkJY14jVMiRk9ysnq1Sz/VZlSOxx+D3M828sxy8dMKuk
dDhwgZmiidlvSx6cnfutIJBqo1dBXy/h0GN3p+wSp9ZdrKpaIZLmrGO2vNOSIN9f/M6qzjocylPA
fW57PCsljpGBnnV77OaMamKOt629Ka45i+Xv+u6EpL1uNzrdUToMwFW7LCEfZQp9XK4HU/MXX3hT
lu+aNvPKPEX3LSql2tB0L1azJGTfdCONW7Ql2WBU95Z/B+wecbAD9VaUjZp1L40tP57eiNCuuCh4
SGelfFzivh9PdiZryzljCI5eBQnkYNX94n3xn4R+rv+JoO3fLLUYLCbKt74iWhux5ZkxAymsChBN
J4g4HeOYQehKjAk49dzX2bVTngFOc2lBkiqTak/y9kgfmzk1QtYalPFjZsh15kUkwpW4cScML6ZU
yuAkXDAFjdXQ1fnvWOqzVMzC7SaHbtDTiu1mkiWe9/imk05M0LBlMsoOwWm3f5tV/qckL4yNS2Q0
PQk2jtGXMCJ4bI7WD+wYYmD0JFn6vWx/BxpMDCDPHbSoqRCeeDQmZm0ioPl663bcuLg1h52Ew9Ua
Vn47D1KNmulfIdPU4Njr3qqieJtoO3SIIZpaaBcQHUvYjIMAVS9FQ55sxJGCeoY6t3M78wGPvmZA
61V2QExpns8+SZgCMeebTmUD9cB1OX2J0sTwk7uZvPCt7oT/WeYV66REYUP7tovOZoc8bvLkcDFI
J3gkg3Pf6Vksqmq3f3cj1X50m+HpEaiqbhTSKVPA6cBUmskgM0YegierXopve16oDC05G/gS7Pqv
TIglxVylD6vwkc1aJseFfH7zQNOvhBe4LxUZ1S+2nwZV9Nvz/LvdmONHGug6x7sKjpWBktg3J6fd
uyWDqKpijWpzVKc+RcTAxFT/krRPSRalGT/aZ6b7zF6zCdKm+UumH9wQXm8B/rNtkNd22Jtjdcdf
OTrzTsYShKzDpP8wBqaIchwncKTXvhFAm/DU1xpllDCDyCtMfUUDI2j8Nqrvzvc/lEBgDUGIoWfb
QSYPcnMMlNxymWecjS6TijtifvPR/zBDDRE3G9uyZQE55/a+e60iMTHptQg9AgkqiI4QsyUjswPg
+lUn+vdd75elU0pv1ZoYSxFVzLX7zLJg11rxHw3dfcAIRRGPpf9eZgWYmoV12dbfZ2DtGF3KHht3
txh3v5MJFRPqk1BjplSdk4s79PySf0kxYjD+Fgr/z46as86omPf8HDNcc6N28INcQiZpP4Ma9Jjl
yDZh+UBY3T3cdglGHBVpPcJ6A4eAIieDiTMXB7ZNh+1p6rEPz7k+TsyNKzgKwxgbtfqeYeLqfY6s
n56/LlhK6p3P6jvaL9SvxtCKJg1juaJJG/B1viiRjMEZJqz1Oe6BxX1jofh1EbF39wkUCctfz93+
lnjdO4wb5sxQQAyOY5z13nsdjgsuCk0W8A4r+VWyI/7WsI7zM2BlnX0z4JQj/DnR+o/LTH9Gkikf
cSR0KnOcEUuJ2udjFT/XVqIU/9XaLwK5jyMCaurXyLw6jAGfH33dGXoO/pESogFNoSG0sOQzMUeW
JTitIONwOBiZAQRLeDAs+W5c/zb23Hl5kKYTa5d3hKLHXZeYk32zMWFLsI2BvvQNxrVKb+O0CkuB
/x6JyzuoqcP3MQUuB/irsubTtzQD3og8VMaUF/uJQFBdksPuo31woQLwTSX0496r4iCeX4iGC5WW
YFSQV4yHUhtEZmh9Fix2SkQYtHJw75zdCyQhaW+52yZEube37CQq4o4XQX3lCVgHA/ExhmXe0f60
Ub5lMt0vraA5hiYktQ5DnjQ8GmueUNys0hpJ05Ou7MXfhzTxCUPRVmNZPsq4aOZVvYX3b5nTfztl
yJ7UGqM6czNdPX0fLWkW/BEysNvPF3MKUY/sNIgoDK9TdDrcJXweYMMcaunXZO2ig8cu2/RRU8aZ
0KUE+zTrbzpKFwmnM4UDWRS1Vhuk+nqLlNLpBIyzIrqyE5DdO+CSzm01Y5TT+ZQWztIkGwmnx2AK
ixNlArRHp+rzp3wUKxcej0UrNUXMa60/dFkAqUHiVGyz9Ll6t2Xg9pju9kYATQwBUwb9rKE0vGR+
5cnFJqOziCD3sgYCr6zGq3DAckaHheHBpRSmWWadjM5eh4F/gXEOqetO5rX6fAVipNt/BesWh5ES
finLd8Qg+R77yGnt4M+nQni8qW68N0UPm73j+FUh0/XMoqOfU1UGRFCEuO+GUer5csNu6QMOXiIM
Aw6BH6gJBhk9/YtdXlCWSprdq/T85lp2FJSVRAkMSrluAYks1KTgGZYGu586H3CY2OVvUKMHS57X
RqiSvlJX6nurR2Il+di04BkKvAHukNIKFwCF/g3MvvU6Xd9IBwxjuNWPH6wMEwLeCJDia9LnRZsc
SI1yGAziV+6stUmipoCxVVYmGV9BvuXEoAnADPGAnC/ecDilo/VkRpECtjaVvZRVx3e2hxOYqaaD
Cn7loRv65qy1NeqYZAn97itScwmy19ojqNT1AqltRmLVL1zdHY0+X7+ewuWX0DmZESG2VRJjRDfu
Hcupq/z4YXOEV5zF4wuUAbSjSLThtmz/2l8/oB1XKLaIELgpkVh2g+mYIZPpZGA2jUQP4fpOQ10n
lM9te+MZaeTSHq4+PqqaBq8SGs5IyWfK9fBdPULZv12OdTDeAeDm9c14liPOKHUjADeqleycKBda
0sG6MoKsEK4HAUvb+aCUwlFNFHus9ZOwPRDdHLBRK+v9Q7Ct4mtKvk01sZaFI5+PykczXOjTHDr3
mnpL25wiwOhu72ek1qpig672vKvKtA4cWoKlMjXn5ZxQWzuj1AsDMLmketFLKjjHxKj7FM6rRP9+
0lfEeIwh0ucE+K5fOGUDgYsPS91zEpHADrObAwPkLhD2LQ1azh1PL+FJ3vmUzqv5RRMcQ2sCqAXI
w69KpQwIs4Uot6SAm1ryG1L+OoQ1mCEmEgPaq+JW6emU7DyoQs3/bCvDKZI9c6CxMtV85RrEcT5+
8wxtELece2Y0qe9jcYvH5AWMqSd77iIgn/VSuf4GExa4VpMmK2JPRVLV0yL66Vb0QpBNPvhDhQfN
ZpTvnFTxFsPNaNXucSFl5DQCtMLD6Z5oKwHNHBEGeIm1vTNZDJnnBRtY/nmxSd42eKFo4maG4cuD
4a83tdV1a6UrpvJhOfR0OVw3v1okOBGbX2W6tvwtVej5wA57vIW30W4EQaXv2cWiRcKY9qsDOCUL
2C4EaNJ8jimZa5xzdX9n0witJxxl/79113b+1sVLpMJj1If3mlDD5ZbqD2dAMBkuLsIY0YQHK0Ci
JBgeBvM2xLzSlieq1QoqSA/kSWRPRBukLYtHaGLqg77EBVuryR5fKu0KPR8aS7/tot0dcpV4zqUA
RU0y9NnMIPjpySsQwmTg7csNCFP0SW30RwTJxK8ZQFIQtC16HOygvI86BzjUPGLUvcfag/u/U06m
neOa0k43KFThOJytUjP7J1VSNxI9ECd2hOqz9LAg2qTdsFZTwteXH2BA3GJyE4qLs+M1DWyJfdza
P1yvEmpKKOFdKXU7bNWgiSOY1DJ/jGrxxTFqYWh0d5LPfVCwPddsBIBPxsD5fAtJhmYqW5Vy5Uv9
HqW4MfKPAROSQ9pwI7G65Ru/Dp4Wg24EKUiR8y38EIUMIa2lJcPZjxL/oZ5HJwJnn/OWAT+habC7
l7IDclHt91jCNCF59ePaATPOxZfcB0Kivp1gteA0bWvk7ubPGWRwtJwAQWinIkM14HuxqAvndXae
Y61zmTBNnh1Dh47azY/EKidLpk4ohfdRxkwmlVG6FVYDp8GvbZSfakzCT6BAId2l7s6dRRqEkLX3
gIy1Y3M+kfdSUbCw/O0b5Lnwy4PJyF9u5eFgsFWL7rHv5/798Wz4Ymlb0qXv3qD5/THGZF88KG0h
2iXSLlMmqI6Ee0n75aMI8mwntLvCAOCiZzgGYt67GQxX4ov/DqYXfmt426MLdmzaf35JH7TK64XN
ObOb1hcvR5Ja2O8hBtDo+/sdre1J75e3qHkFQBdHKRFa2I1PtpiTyds0/LIUM+xJjFSumVS+yJ2M
7Ilw0tyTPpDGk2xn0FrmqHE2/9Rmgcjanah8OJ6JxDtw98NWwLgyyrPL4G/BCxxndszXlm+Emnyg
INp/eE7+0ToNojMv9uMfUdujasAU1F6SA1Bwtbm6E4/qrK2QOEItJZeWaDdgShhdAMH6IL54JO4R
rphKno+EZiyRujGc+GE8ev6tSi2HoBXAKq720Xa8hDGd9wt7/HrcqaVIbOliszIBaXtzpVak43mG
Zkp++t2x59SRF+xvQ4Jn3roG2hotWkIy+rQlxzgTwOG4pfvKQd9jOi/+KWwRHIG5F7iXH3i+0wIG
WlcM47gBZjvpfYKC9lma0s5PXjTW868Xs+4UAc+tjJDUTVG7PmAcSLp3aorba1X64vNxFB9lwCYp
+iilGtxgqB8dXrx30OlHK1MGKc/dK9PvKck4k6Y0wrYvnvCPyEo10mp9Gpo5xZiE/M0J9b+1MnTR
FW0blvFMajXtXKZiLg73vppTQbLVKGAHb3gVwWHJtMI+vCsT9O7gBrqkuVhzPp94M4rP64t6vPYf
NqZPeH4jOaZiD+EJCZ72eaNhEUXvKSBg+WUG0mX9cOPiaZKMF9OCt0feJwaS+s/skMamoxLJNZjE
RX4j6xaoiqS5OMjDPp79NuzngG64BhwlYUtr4sxiCvohW5JlOi9tdUuA3iVKNqK6v2QffpD1oAWM
Zl0mlPyZyspXE0GNSBlPmrJBCrxrMARevoAGAuuBSbaFLnnPIFW8ELaNsvp9Fy03SZs8t5wxU350
Dktg1uPsrv0eM1qtnQEiOq5K3ACzlP6DIA9LtYEPsKZDZRfD9rVH5MhlhxrlSpbQYSuECf7f5PI/
Xr6vNlUM0L77Ht/IJeiEOwMeuKKaB+7V9RqiHMim/8hErapGdY1+9E+DLZNjlH4H8q+eIV8U6lAu
j97HFssrW/brb50+q9DlkI36VamtI/8hmdfRl+AcskqIX1IfwHK/ngvfD8ZZ42pfnR5VaL+Awq7g
cc725ByC9sRpeZTxrraahAXhobULvjUu9lMB20RsnMPPQ8NBZtjsWf3A027LiHp6LfYWIf3EYWUN
vsvaaXQePXJ4eRWQmgyNsEiP2yV1ilmNNslLoEXZ/s1HaWuYysQgfcQoIbugUg5fhNJVd+d+p2rt
JJB0zUTyp0CgOqkU6vaIbkPZgnUeRVyQTZuKZEZMOTzmoaEceiD+zDJPYUVgryneLVpG0xvZ7cv7
T6rD0Q7bTBHr5N4yr3M/zQ+rc+C/ep5P+5OTp6yI6tvrDCCxziJRjHynZD+dKif7nglFkYOwA/Lk
9CPIwxnnww2pgwQ9AhiXwOaiCBDB745QaXfcD3hhIjqYRowLoytpRiuokMduknhizMLCvuxsZt+8
IrWXQd8qdXpsysew7Uh7RsQNYXFsDC6yBGYTBJ1cJj97XqhGHiAN8EVRsgpvrHDV9zZkZKZwmd1l
eg1xMxQNwrrFPuVvWhk4k7IG3WHhGdt1yTiKmGqSdkzMwIXgyy9wCQvuIw7sFD0SxOLQjMLEeTZl
feZED+YfC13GR2vQTEJzVlhhF2XJgqaNnGBugwkUl3lKw38PVTQNBtpcSPJw3QONeP/JqINZ4ia9
3gibKFFHqgTK93aL4CYUC9VRjla1j0pMr3OK5/P7hSDI0N/5+URbyVq5U0Jj4EScQJ7AH49p+inF
BxnvniYss2w04lfQNulHktqrDBfVeCMRWGv8aA1IwAwfIXT2ELv6YU0hf59S5IMYGQJOAhF6kaTo
lAlw2D9yjc9FFMthEV0I9r+W4wMFxEw5b3Zw2zFunrUR5+Aryz/D8FltA0cx3XKbbykuhgz2916R
i6ExHrN+5Ulaxai9htR6+ELkxhHGfnZr0+vhzV/DM7AgBWChgSGZfWkP0xTml+u6xSz9zg03jV/Q
p1Y9l3zN647tiZoPmzxnjWtcWssYp1HIWPE7EI6fO7NHlyzRRSmJ76Zh9kTkfnhNKs8xaic2jZ2Z
OVCm7SGWwyEvfxxBmM2bcVZJeLNPHFf3LVEMB0mRElT+CffMtHCbqQ4rOi5G0nNKug03QTtOZiBO
cvkRJKv7MwFndA0CT5Ji5+U9qZVkJ1PRZ8dJUVcGg6bMM0hcuFHj/aA5QTXoEJZrY5dXWvbcL4fX
CqeDk5WDnnOifmzHdbZhV1x+MqGPvWkYWMbjGRKzDAHIoy2rppKkBeySq5tyaxdQC0lWovpklGne
y5crX4K6eo3mbJh9XiIu+TQqbvzbhnlqKs1RK2LYSf4O5D/zOgXbzbQyN80WZjFIRPzw005WPMHE
10b1FxgFc6/GuFfIpVxxW5nfEgslMmBvENGoEnWIn86rxGuBtgLhfY3sIv1OBu5TZq5hkgiKYj3c
gQQ9MvyK/KFO6Ekfs1PCQMQuzUH0Dki8/p+qGR3EJTu05Tq/NRkkQUXsKQ9iQMnuMbLwMkIYLgyN
tghH1SjhJlCXJq1wIwJ3DD/kLzDDfur3Y8QpRYDImOTbLRMbEq1AHJixezKvNb6C9uZMrBItnltd
rrd2C6+xgbHP5t4ySvPjrM/4A8HQNVzJaov7t8hkOe14XDu+quUpByvTXJqLpB6xxF6HPfxaweCW
76+aJTcLZqdd+JXpNxN7uN3+8Xpi3jH3hcpT24cdhClqYdTHrENENGhSdWZy2oB2v6uwDu2TaOOX
ExWwqjVYPfbUT2Z2sQwjSfudGOXT3tAYy0vBI26PcMvWcNT/1JEkRSXEr8cWwuOuKtUqOoR0OXgD
dt/QrcWQSzFctTdLUA7m5iRKv6I3lOvxXcS5WkS6gEu8YxzWiMs4N6ISr5InkWNHtXgWCr3khlUr
dt4rUwGN8MzRqnQnHLmYxOUq1HEuGh7Hh46jlMXmfSzzaopYoBaLKp/vbtUtb81CMJx87FalppwK
T8q3odv1Fc3dabWNfjdypGxdCWmTjbNV0xvnroSHc0Ru2ZbfZ3x7NYpHiEVVmW3aSHFzJdPK4+JW
Vsq/GN2n/+d09lAr3+lN7trVRYI9TkGdYK8iSdqM0v6nBEj3ojnsBo4It45wteKFi4tdYH0GvDDa
S+tNnsO3dcMVE9s/0RWaSWVlOd6b8HY2fr+45LZbGhpe07kw5v1XFCS749ftBtDJfOvC3ImgKhRr
lrHxKddCORgGZsDUz3G3Ebz+Ex51B+8UT3Xjt1CIdzmp4yUZAigM30IqON0qyY34bJ1OJFKe1xBb
npTOfjmQ7Sb6nghPITtqjS/RaR6Qah3sURv79f/DAIZsdSXcLqONarh3hBHi+FmkipzD9QJGyrxX
dE/m2KA5gJ5iqeMUrW+XPak64QcfQizWVWGowaWpTH3W4QBiuHQ5oGcPVGjkrsQBe167Z3jEH0LO
cYyBVzv8zfecZLJfO+lGQq/Lle6dYEgbLQkAwsNUYS58JrZy7WktBQHgjcG27z8eCkRI9AOmj9lW
tLfs+zRLeDTXUs3FO5dH54OFo4PexiTugNeaim+O1GPgjp2NK5VqBdlcjXgPAu5FHaqkfMW/5eBy
qbE268R42eucvvSy34hpaWyOqT16nw+8Cuf2O8OxbyzttY5xOUu0E8EMpJV/vIJtgxTjPdMZPOVF
tKDRXe5qc/gtwa5CqRPLAaSUN7vQOL+0/uHhKC6TAyAZ/GNXR2bUX8bLHFvi7rO81fVmL9A7ItoK
koivbvJAWjbFau4WlOy+HsOovwZ5SU2bvr1w5Pphp7hoNbr/vKMLCLoC7ntvU2bn5dRts+5+ci7F
Trxn/GRD+cEM+k79ylx20hUr5yOVhpVGuTgCub31vzY+qZSjqxgyg/fn3N4ucoN3vtFlZTEHrgN+
yrrhnK/uFjZBZ8hSX2sZtUva3Fzyul29lc/BfbsFwYuFJv8toqf/onTZmmrTiudWUuyZ5VaCY0ow
ikMUMSqXjRhjW+tyS34TLzE+v8sHStNkokExcDiK8MAFSOjoBuwd1cwLf5O7xTedaz4OPf0rTk7P
KnURslcxcK9nccs2Nr+rBsrQEPJbEby249R4Gvseos4qp6ua1J1n/IlOa+FO2M+rjh3eHtm3upZO
26+6eMEvtovwjyTSjnNRGCLhOBy/XcmCwwKBt7iVbpwchFhMwShRPjKS3GMd55OQhxL/3aRbaMtF
5ZAjcMYLZON4iRCyJbsTyNwdraEKWgkdpExKT8JQcmDfLbjVQCbrbZXSKWks2+tKR3YzV9vhNCT2
1P0Yv6ZwAO1+wL0HK0aCWwBfYTsvitZP8qbKshDCsESxcOFQtWG5VvszGSuzddMcu3Q84UTStJY7
ZPkaQ5s1gXUAczWXCwjyHsP3vT9J4pilvYwEscQnMHUEEekRb7u9hVJcshS+pEUVhoInpCdYpY8d
/d68QM6roXZaGrS3J0+aYLXsbHJ36Yl3eX8goYBxWU10LH+fGUbAq3BdL000w5vYTkp2x0buKVqR
9Kq8DvFmMmG5W+StjHSy+nbpq79xelMPDvrS7z8J1q1R6nkS7yY0iS1pW2okFNf1mXvLm6SRMcAi
zhwYvERzOmondT00FTSN5s3LCMw8klEhXYEPhf6l+OI9tNMNzLoZROC1kcYPstHsSdySfFOl1m4y
DQJFuuja97k9RTfMISOc5eMwdwtnwrrVz2+V7zQG1rsA69w2FKptyvjHaAMNXN+dsl31+vcQOui9
CxwfAOO0mpo9OKzKPGs1NdnalpQbAXmsV7wnFeJBACCVmLU9PJqT3iCxxywN0dsnoxnQ+nxadYBZ
es5w8gKjEfGRdPrU60uUiEpknLLsVXQhi4qG33qkmdN0jyL3oocDW2NW9oEPku0X/TtbwB8CIaEa
R7ZOz0alhTjAyaQh0Gk5KTdzNCbEF/Ctd9qZCuOFHdQy3gFWl+TBqP7RTq/6oQ8j8X8voprDOLiC
9ODTo1vE0QCFZfMmb1TWVX5efvLU0SeXxAXsqJH6QsO2ePEOrH1wO3ziJM0CJgV6C/AQoPmB43RT
3Koec2+7cZBQt1TMxXGigy+rekv7WnGTV/EK5itXEnvVhuDb1ZpP9qnMyIupMph0I0o985UxZ1yE
ZoQfRJ+Sf7wIGd1/vZClINTsYHQBpBclAAw4+XzZSsAfJncW2lwxAgAbg9HUHj4wW8nKCs/y0i7x
G5SpwoR22zHrCuYAZ2hr5FQlNhnYmWilIc8FNtQRPwxOtWR/ekSwPT1gDiVR+/KQWpaKKeqR6Cop
TcL9n+Nkd9nfSmvXH1f41V5LYEJJIUiIBbYtOqf9ShgqPmwhnDJVwfUT1PaI4G4GfNvZgPCpLIaO
SlAZSZkbMRN7gRoITn4SqeAAC+BLRNhE6weiAs4TQe4vpdP2cH/a4m3ivVP2Xjhr+9VGpQxk2we5
xpvp1qne1IVSJvFBe4NYArle4eMtYRDKl2nzz/7IihGmDFWnrl4h5Wl7ReGpaZZK6cxjRW/S5o7J
ZD7D5hHqFDJtJ3BEbC1qBBa7WBCOwkrC+/IOc0LOMCprCjCXPpDliRNAM8w25xDp/tYQRRsemAQg
Tkx2H/kMYzZJMw51iXiLXMtAL4VXNQOHtsNRsVFbRthuXAbxPWcgz2IA37TeBmnbqe2N/BbAeqM3
Uek+xQRXkCPnh4DeZLFt9n9r22AE/vKoyxgniLoqlFYjutPhdOjajSRkMQGU81BMynf72Wy7Nz9f
bzeD3V5JOrW0ICLHuF4+jAvSW/Ahj5/R9X4YeNpSxy5HyxnaBOnjrOhqGCzfC8m6wEMDU+K8Dn2Z
I/UMCmE4N0cAqIKOitKhGNdgTzMPto1xwATiI9AwfrFb3PA2SCetuor7BbAlt1pU0TaUIlsvBz5I
12qxylafuJtNDCAcuNbueNaSB+Q+w43PUBcPRWjfUyI8Q8uI3tJkhzZsLsDwqeAt1662uTvWtEL4
GN7XGEpf0Ceptbw2Zvgm+PTqvbyas2e+lAjOTcko0gyxkvoDXc03N7faaoth+9RZtY3uXLjw5Dor
wsZrrlBUwVKFFMlxWHOcNq51gI1O/bSvMT4aVKZEY+e2seFxmfAmbI3gAvBqSvPWAHzb4Jg7+3CL
r4TtEIEBCrU5LaF8FCwxZoG7tFoYYEu/HL6OHZ/RPdEZ/TEot44WRMnIwpm6G89DomwpLMbF5ZGr
mGbqd5jyiWxLOS79pKAhP1FapaNvaijcV72gAlm1emLJBzOn4NRtSwzleqKdMdU/oQ8C4o9BNbwB
76M2ZpOVci/ZiYJeQqVl4c6HE9DjAlaiOJn7hUoucayiRbLE3b2ZdOoZaZmZFdnpzu+G50OW7PHG
dix+PirSp5sgXJLPwdCh5lc4v1woTsRbGZegmh4FTW8k3OvyCDjapS3idOvc0NnPB+v16i/nLmuT
asXdONAqaBXK1F+YLku3IrO4HoPvBhRhr+LUwwB3YRmLZgdK19U79ToTHr4qYiGqBU3SkjxM8Vnu
qvYHeDTa8V1RPfFeAxlwnQFZ+xaFBNIAxMPgfDhbvm0b25dzV6r7IoKhuhz1miQCpxKNS095jaIt
1sTRzNf+FgHUfiVJTYDIUOE148tJM8uzsFyeP+ZBLGg4FRHvevACDAG6Y4PACL4v8N2plcjgN+2e
4ABuNnh2HVFPcc/BmUD50FTwKFvVOf1o8nZSnj0mblrXab2xrWH40f/bSqRzpUm9g2zO49yCnoXA
p3+upQwYmavhW11OjsCkBEEAfuaekhuTMiLIjfsgUoBGK3pveHky0EyGdbHKaz6MDkYxmHoLF1Zu
tlvuzjwmzL5i+BZ+xDElVYnCEm1KNw8fuyXsXiHy4GWmaz3Pb99gM0dAqMyShn8B/uQVBWK6mgGb
QYThc+m4WcGjof277tJXyxzjpk//uNrfjzQDZTT4mWCjcTxE9YyoIsHyO+knPDoQ34+erPGya0yD
sJcbGaiCngOX9OBTi1MkKWOiMj9vcC4FvXnWFiiDRHxTKTGJJ1lbWChcaXmo0E/9eXjliFwYdFWO
tnQkhGhl7Jo2oy3o/PpLtWK92/dVzyslkyBTSVI7DJKXoA92F9LHSq0MZirQPguUEx4CwNOq39lj
IdypR8fgWjWThKAyxmlFtYDvm4IVEDjX/uNKdnsRbhIlRKLUNFMyht2G2Qzr2N1ELWGTs4AT8MMb
bprFlw3pHqjNTjBRPYksBrrU9j1HjJoEx9HqaTIa6gm112RkWqDAqgJruVQj0zgjNeyS6bT/sqW1
T6jdVZjcdUUOZkQsL20uzO8ZetrjcBQ01PL/29PqWh3d3s06P6zuzIArj0C1FRRDcsmeeC/GaKQx
CkMdJsvoKenaq2cZSw15H/KcFkNAZEGW7u8ieB/bG3XIQdt9wRYgrtrCnB2xR3Kq6vDfWxT0ecuN
zsqBBOB64QfR729ePcaAFMYi2907X6TCcmqmJZVPaoP9vuewsgW2uOYCIzFDbNaEulb+xhj1A0DP
apOqaw0KUHKoY+DXmgp26l7LVGKOS4KZdzLIf764x+NDmTjbYq/PcirJ5Hmc+YViEOsfyvm7jJtc
QgisNT35ZDF9BV5LQJoj2Xyhj7iHfQUFcizAL/8FXLmXIJSh18gGsLsogqdPDbDpmhq6HRAmXhJV
88BSFxCxY1WbZhaxpJvNhyVVWD0UA3dq97b93cisuf6o+OmYGkeBmGfbFqz9f1f9uSVruwReCJKu
xV2V7UmZSLY8HUUtOWXF5hHUURU4DUZd4tfozYGpM1fGy9/o2WTmGzwCO4e3UsZJLYI+L9JHKjdW
vjrJR4tJ+XUfe5bU1hbHcFfYFgJ0NW/tOBqTyIe7WS7EPS/HEsodBJnlKOFXMQMzo10BeFOAbK8L
hxPOOsc23nxcQEbkNYXNtREUeEpCFM56A7MzIBSSX0So9pchkGbmpgOppzFDgyrt6BlgQ6m0Z6As
tTpscvq7VI/pFUWcIsOzZjQCTb9rM/zG2193XN2yezf1jXyvu4JyuMySkanvh0EJCZWyhpOg5+XL
83YqPhALt0YipGy8E1hWpzxSaQF8BNbDIVrXHJ3WwN2JkrOhTdrH39zquJuNLXJXlK/deBGT4b8A
yQveC/PZDIxANZAlCOVzRqOY2FxyPLWuEC6Zl73rgn7/ciP3CqB19tUXPhKV/BcZ9t5g3b0Ey2LJ
nCKNr4HeZyWSosJCm0aJFxNiNDBcghxTd0hVme45oLLYZUa0aVUktv+iecFAt/BPd4MmZQAxsPKP
GZhJyxDa55kIyMqLpP9CYP2Ne86ql2jMWQqiSO+zeF9sTyfnJb/nc00bJaU12w1zWgxX4vNXSzV4
5Shq0puIfdMGDpv/S+JrYTOCoqwhlgy2FLETahGtPGL1K4nDDe5SQEIwhqtUGDi9ttV0cJBOkCU8
HRJZZV7RJb/63eMDJBZYBm8Q4ZQ/gnw1QJ/102SzzdCVs0NTbs9Iw+vfQj8TS12Xd0CqncxiIg+G
T1DroSfODXCWJ8egB7+H3zyXuIyxKp/pmU6+Mp08aJiGmHd6hZALWkK+vemV8aZtayh6bHsk9K16
VeTipcvYKjK6uIokChyF4FwKKq6kBWvL7gqMKRpSvhdQreFRz8U3NKIDGots5X7tGDf1wuj5j4hY
1217NwCedvXdbsuNXvACXjZhQRDuT44qIHgdKyDmS1pTfBsk3M9Pt/iZ3NeafD56dCIq6mgYtEFX
XZiUqdNLreKTpnsMIXZ62xFhrWD7TvkLY6uxKL0ctWSMA7ntNcTncPe3k+IJ3CJS+4f0cqWdCE2m
gG9hzlK5DhbpXBPs+N+sRj2lfolNx/C74rcUmF/NxdHFcYkSi9PMJO90qMFAhFFu884cDHil7eLa
9Tl4ziiczmJAjW3wMY9JNpS46qRtQuPsaY4DXc0oWUkhCFZ/0e/wXxgXfHuuXEEZ1bJMvIFlUO6c
ILfvZOPN7a0U9UcrNS9BP0+kytM0d1WVJ6uJ3wnBtvXLdKqo5X4Wail12bCE40euz7PZAUdimrKn
jjzzTvav2Uqy1k66Bkp6LoabiLFHr+p5ZtLwPuoMwN0kiaR/OdG2CU1ApZ0lRbXrazdEFRZ6iyvh
QM9BRV7nLtveVowMFJzQFHrpUOk1bnxWQ7qF1p/+jhWsHmEwCA8DQZpA8wAGIzrZjaBqoRKBgloJ
H6RFXSbwW/HKPknKMu69I8cOYfPLcoyWpYezOx5d247hKvLvI2WLVTlCIR2ilOlEZgkEvtNMaaPN
7ozhPqEgEfGr9ISCqPUlGuDsiyHQya0hGmMGZXGUbrUlyn5DqI79Qv/yHzwM08Qd9vlG4m33XUR9
CzlqLR+jQynbAWTNpHcRHy+qRkCdvATJqpO8Zv6lw5vtOhkGsDCJhENY0yFYT2VJYH2rAI/HSzd6
ZF0BB6gFKZN9KF168SE917LDvgvfvay4xm/qSdXdPE5QMNgICBpTIknsdHuEso8agTEdbVo0n8fd
7cGqdYUTiJa6BqqrFZz/WHFYA72XBmUUyPSrKSKnMwmp5pQvQkCdNmqxpllbEF90Lf6/AGY7wDwT
cd9YNjQ8udi+IQ7WivHJKE+whqk6HpcKR1tdGrQL3B+GGu2RE/34uLHHxZoOiXFg/F5YVCyDgxss
n5FjTHd0x7286934QVCavsz3fdkcuBxwO8k01owj2U+3oQLvaIITj25zPaMr6x+af50f5M15pq3S
vjAW30wqkP6S0/NqC42jXpZGdiLVU/XpxpMYXh8rSYMWDvu9AjUZ0z7LX/TY7WdXrBUc8S2BdEhj
8FEDQwCO9snQTJphapb+JGIHGqYgvVCK/5gHdP8PtW1KyW1QtV8Mg7Q6ZmbgiWdzwlC4h1S7Eikp
5sACkKVfkKAPfCz7pG/0u+zYUIesbRJL5ifPg7iFHZxIlo2IYXAu8t/Z9PMkEwp5qSnF+cQ87scl
aZAlfCHI8rJbUaoFeSskENv3NEB+0AfiL08r69Wm5c/VwH7iMOV7PiHKtE0XjdQ/NihEDxQRzuNG
dcgwvI9W1Cx09SoS1zLaFp7gEFCBhtfPVyjAwzuGr5EBuzwWOSTCy7QYSf72pfKj4JWZbD0fcTHx
lP41R76+VF7y4x9VfH5z8H8oyV2wSuceCGJB04RObIad2nR/wA2NIJ8+5vF3C1Y8tT+kL7DKKjVw
b2J8V+DjBE3ezZopfs2jq/3qLIPR/xThA7LmCc+MHAVAvg4aLBhQ8ccd3uFCFA2oqKnwofVamBdK
VUcRAZnTz1mLy8EBuqjSfULsD5JC6bCWb+iqj9ykZQe+ZZgfMcZjAslKorg8ZahkPE6yulpnZmsp
ZDuz8sfqhUmAz+p/7ApDfT8uPOrgTWkcRy1KC56Rs8uSmb9dONPsfySUgY9DgROkvbfNCSHviGSN
2PbdEyHAbw++htvhNCP27F8Ojd7QFxuFofKQFHT1tpO8uAXoG5zWFaGo5xZXpzI0tFbs9nPsm3n4
DZoe22u40THZbksJHo+WzEKakHYJm9NOht5ooH/MjccwUruD/YXRvxry325GjV96YoAaYrRxY9DL
fP7O2xkte4ElISgITX1s//N+UgLru3vngWf+I9UEa44cRQY71jKE1ZtIInwdEpAoStWzx4sPwffl
hGEo8Iq0XI5tqMHjc972UcUZAu95hgQkVjHXI5RISV2Uihat9W9/R/M0HpQzSW9LcVCUuUbznIH1
6uTOBzxx46yJjDmFOJiKPgw+ryB6YW/vtuQvnW7Jb+RoJme56ot8uR4Swp4XXg4AG55ohH22EKW6
w4T2eQdY24WjzSHZ4b6osAK/rIFtT1RS5YaboXjV6M+hrU7sVyw2/+zqNcXk0eFi22KKu/vLCFg1
6VM4Kgm7NTpgX6yGOwta6mA868VuXTM5Za7YOYRLvxhZzZJP2VJredJlCZN8Yb5NAce6biiW/Pkj
4KJbVq6GfDp8CCH6BuIDZNGYUI1ipWnj9Modb42vLU5huplQRn5Ud1WEgATSpEOtltWl52atgf68
Anl0FC0s+IAyoevNRGf4gSmnjnSq1KCTNZ7HlB/cea2HK+9CPX8YsezIKcSYUNhtXjPPaaWRbMMe
A1JQo2u2v3B03qsO68EiF9KNwzgur8mVd/JQQU9f8vInJoPUd5kxCmZhDOXIps4zQiXBdfyYps8d
4/NoK2zAiGPCTASn5t6MNpwJuYgPwSNMP8ClqJz/Jf6AYTanikq9UFacqxzo//pa0RYGfiuO05or
/Km3QS0SczWcg4zFKP4xPOATsAgygjlI1gHjbWiprafjO2pD/7rdmr8/OINt9Uoq0HE0gIRBv7Qx
2ofOar6jPF2Gll0e1HcFD1xQmgDrGASj9QQz9kToGTvJTYs2+gY81Z8SypzQQxm2Ag1X99pV88g8
RYVElwLfcjE9gY+m6KG3kiWGE4I9RxB8hVRrR6BK5PBI1ycfs1f8uikeGjBPuKXl8+OZwuIyehtP
Kr/TdfyGcQKy2KaUsDARdwIP0T35PwBVW8qKUjRTuqDg5Sz4TSwyig4eHfga5Xvn4IdYMVigGtts
XQ1gBpcWVEP2sxVr+fMxKlToe1b2+mrtNPvOcKK2Pc/w3S30Mo4g7Ozj3KhhMs3OMuXxKcaHNavC
6v19J6eQNtwfcftTOVIMjr7j3PQNj8xAjKcyjQxARI2hD8y//+Uc75XTcyuuZWcgt12uuvOjwNbI
IlWFjrqN8SBaKb4synKhTfO1WluCeYl2BGSHFWRHk09iEes2y3P2KUTW8yW+32URxWL8WtHF54PV
uEdnDr2O2FbqQoCJB86JK9GVcgm69pN3wuzYUROSxIiFu5XgFcM1aGcjzeEZDveamu4JwPon/ayE
WnN/sMks6vvaZNhHd7Kr9HGcfXJmJWAX2OlOWv/t2R2KwNMYzpkAIuamiEgzTI8HLdnDll3gVpVQ
jo9NkpzSXMe0aU3MVSr+Mh1QW5XDrkKBOYMGOBqINOSL28nNBy8D2lyMBbnuVtDXVTU2lV6IubJe
K9S7XPX1EtOMBuEegLD0FHMl+mncfzliDCFSWX4Aa8KbF0k/th8fXDM5h9YN5e4LO5NI+LyBVD68
uu0FG2Q3jKwKY6Uu5BqCFWMRi/61O1/eAnQ5ti30cmvpcXzlF2qpU4YlLpXRxlenh0F5MLXgDiWv
p7PrvVgdMx2OnlkIqIlVgOyt7gAAYACdeFKEEKLtLSOpEaMMkf4ADnPPc8+Awrqs81ACZT/uuWoj
hncMj17/DqoLvt8eE//fwUu46AHHHpRcHwp7g7HKFq31Dkl+Sihisn32AvsdU2AWAASAaGG5O2Mj
WGvVQNiime59mwIds1TeZZ5ddP+mn+Etrk1bd9olhEftq3GOrH782pa6C5oSzJZWiH1swHeT1ux+
vo7nOLcw51PzjLFPryjRa5x9FVOnr1tsdlYGM1Bvj7kFnyW+57a49c6XQ0vZTR3hRk4TnUmuq8Bg
fO9IIpg207NaQNj34yOdQ6vKs1vF26ZBN0nv2dZQQVdzmfWuVfWt7Cin6mj3LRGN1k5v8zLF1j8C
4gwv58c1ITnArUC43WKL8enEnY162m4dc77sF1z17Hr+3M5r3Us7cFlm7/niXXvKSR3StejZP8Wb
MVA3P10cEE/C8KK4REExIdCl6EkUJGtL6EU23z6+wzpRCgl7fMr4HZWxr8SFCeBdSTskjXIH5z1Z
Jzm0mhcEuRpcrUeDtE0wLG3wiA43/v9TYRhppYBxa/AWwk+voomiyjKyC02qpc+Uht04sevjhfTb
8hR0VzMdtpE8P8W9lOVLrAvlYvLglELB4aRFzQUNLnp5+CjtVR2MthpBZeFbic5I6ACNdTAd05WJ
QUGX9B78oxDrRlcD61Wum3bTXcdz5YrwYEkzJ0ZHQg6G0gzj0zijBunJEOgomuB6YfXDdyHzDdQ0
grtTb0YvSEtam7VjnFSKixmKgSGOuaaMIjA+rzU56PDOKwuFg4LH+gv2JKWbUKbE8zOUnZbB25zv
643z/IrHDtXkx9WjoMB+PSbDJOlLj4lLagOUrWrMZgrIt33E/tpQL5uUqgH4kHOF4MLQK/Tpk7NN
uIoOXwNmhccE/SxHjFMpKtqXb1JGiy67vcsba0ZuTHZLXs5TCEBKIS/jPHhmf1gFbErQLB6QyTni
mLm+AleFyEPr309Hl2K1M3z8o/2i1Wl2e7a4kKhqB4I/C1fGlqPC7HaKC5FYgXcWWlHRXatTpvOO
A/inqlHjh9v/t+b3eIrHFieFUkmC7+mzBoh1FPcCtZXsesDF7DSVFROrlcwHrDQn/Z4qSjQX2n5G
yeK7wmPYEbfQmAGdHpn8EvI1x5hy05DKjcpi3c452VCCBE5QBQiUITCS7UUs90+6NEqch6ipmAYG
T/eQ+JrOwOBnw+w4RPx89HX3Fo9FzAli5USqdmGC6Z50oc4RD/Tj1zRmj7hbeCNioJXfQ2yjpuYB
tQOKLiO8heVWcYLKs2gS2VfMhSjvydq14uc8cQWv3DyJY7HNkMnNLidQ7Q1LEQEyKKDTesPjtjQp
4UpAiKrI+kazSJIeQeCyN9fnFjZLBtYunpQGoraDoo03qhzahXVJsrAqE/U/1W/5BwbyR5gHFJMH
PMDFS/5UIiIPubazgpR4EwRSbNfpzzwe2vFOP2M4fh9I3Be7l7lJD4ds3vLUERS7e5f+YWLVSlJh
1kJMQdKRw1UwtEQ0uIrTOhLH2HwSOdb6NN+AAo7LblTt+CZfUvucRynn58ATecokUl32uIsex961
UX69WQjTVvmFpu+V+Pa/6mzreqZIXb0JXPGiSsdnNRRLQod30ZdIMWJRsd1Tq3mGzr5fAoG9B1aH
KzfFma8EK8A3GVnu4kTOSdSBDuYdse1Jz46KcYohsTRZXeItK4UoYwKEEqtwNLxMWf2iKx7Tn4Xf
2lmMlOHxQe+LO91QXffyfPsWVQx2TBoR/p3y8wD1BDcdvzo4gJyS9t7lwDZ8A21hj0HuL5tAit8l
SzDDtt93zCTi7lhGJz66bX0T2TFzHawwaUUGObgaoSTq3XmdI97Lv5jccO4t5jbeaFJyMLhSLUMH
uVtVDCpLCxnhFcB2Ep9KFzZt45CvD/FeI3Srx+QcArtNjPnG8xqkV08JAYxani3IZHjfZiZofKuO
YH/zayrx2YJR0zgCwQREXKd6SmAzjlMg/wq1g+aGlehQvIea+lJrFiP1dz/qcDIJx15rYkzvl6h+
d/goXVZnrB9k+xdBd5+1o8ZP4vwIVqp0e5IpWcZ9t59CwCFFLKFFoa4XOMve78LaWLzDwfGSbCLK
xWFQEF9eb+lppLyVqzqf9q7nA9LvTDj3AoEHXRvZsXybhTN+Tx/LPOKLtgLj1UUYGgV8/YVnkJO+
YkskZWePBGD723PtQsu+S85Gsp76CMB3n7H1w8nF1aAtVJwc+bQ0KTbcqwJ9tZr8gXwja207Xx7/
hi/hUeAMxw79NGYdwGKiO/NFv/sBoQPMginDzTwdPNtSVHabEM9lJErdoPVBDAsziNkr4Xb+1O7T
pVVKpXokkcyYP4swxVngEwKnUlsFOhsGPShXr++UfMaAxwl9MwPDveptZxKijIlELejJ7+R+JUm3
SDSNKl9Nh2Mn+M1w6nagOJqnHfiaIMCitVUFye4uaDWkZBtgcPBwO5LalTtINUbP2826PgBHIfk2
M2HZ1Bu1/iM7ZZHkSQ0KbdbrWCc5xSO9kWv/EvfbvqP7GclqKrzORWX63SDELdDrCr9fxsw46w59
GqYDj5nbFK8bl/+pvl5DS9aWP5Oi3Tcehem0MNWzdWFAPfyi1mD/uABD1o1QFx12704a50Og3T5v
h7UARwSAcIxNKcSXDZ2cKPLQIyIAjqo806LSCseR0IkTJN2mMuOb6H8rgQ6Du7Sw7WlqWpsy1G2I
PCvS0fXG09j2IG9wzgxzZJS4D9IiZtpwPdtvHk8qXUVDfA2LTTAWU5HVp9ojoztWSUawC7gCvIhF
OuXSwk9u9AdQFg/Y8nTMSPymiUaTb1Aa/5IZXXJD4VYET3zgkYlC/He+fDT0YhNYr3DYH4khb6Jd
cfUEc9qJZdwHwgC2Hc06HxtY/6xkaAkd9uEBUpaDOFHOLIKPV4jb4iACz1HaKzhYQTqfyq9dixu/
ZOP3x+aQG+t6uZk3PFzTTNEW+H92HaBT3HAJrCZ69bVpDo+GKuH+Xj2ntpMXkW8FE8lfg9WQtga0
2XqmTCg1MUtmHubHEyb5OnZ9FOp7uN+YU+7rEKCa8pMXHnXnXH79U2hel7LnvqUpTpZzPw2aBIlk
xI/C+KPeWgPEWxJNEjCtH5E/6x2TnbyquYC1Bcl4M6y/e7jzibsFye/x0NvWotA7OoKO6q6PkWyy
Iv/cARC462U3XAkHYWQJZSADdZ3k9dxWm2Z+QRmVj++9huluAVFcdpTkXKlX9lzbQYmO4Mnrapk8
9sQMhIdLgQVPgSk2V33T5ibw6QDBmWHc2ngcTiR01DvsOvkUr8C3GXyc6CxVDL+2uZD91gHOrl7T
1VIyXd9BHA523jvAwoHVmKyQpeyu+khprSVtaG6GiGInY5Ls4Fw1mIiVIHFbuxRfOJgthLvwNeCP
31XqLY5YZCvCWCR5ovCtO2i3ac81g/XZp34tSwZN9F89rCEsYYE5KLJnrV3MMJFhgGT7aE0sS2Dy
/uq5N/p7nBsLEQj5tUPLHPVbgfVnZvRMFflv+wCFdcnkq2q7VXJOXEbfkNDA40parSDKNOlDlVZ/
4+dY3DkzNpmU1ogXW8YjUqaV/enFZgmqHJpBph1awhyeYuf65qkx0kymrQ9+qhZdTlfmUEZBMnS2
PxBWRFfWCyByU79HgYLpg/fz3jYXCDM1m1gBpZ+PZelz3JBptFQQ0wBr9LCjvwwNO70jMJ1BsztN
AHXAi3goR52lG/2fzhvP3G3NIUAaSWsd5FDn5hwS5qOpqQkKt9dbaQsPWDVus6RksTyygB/iPfB1
xkjx+iRBYmYvQpPOEXm23NUlmJDlNlJgS7AMztxDkAIsv1UTJuFDOdm//W4qnwBrwMv955AoNQb9
tXAPBBH8o18A3RGAqUhYpWrRehgIt+cDjQmkmaPcE8O8UmZ9IiVfK+DhmZSNyNRSb2e10103twj2
/rhfZPcifaa4jqFwM+96ZO5xFt0rOgkHELKSp1Dvz64irjLnjaYRJFp0eNBL/+r6iODux8w7X6EA
4tMXchnt9YU5xCSygn/5JJMJy2fgY7iSPeQR7USaWtAW53FyR+ZyO9rUshB6PPNH/KM0fhRfotJQ
gWywU2ts+cmElhWkAngwcFnEfgoeLbdpw2FnAi5AMiQilpWkSmQm28RWbaHa/4avi6i+6W1TPFcm
M3MKTUbwkpVejTc1Kvsr6Cl5IAVV53oxAuY30zqRCKn6/tm99Qb6xU04CoeQvVYElBBZWP0X5ES5
6Xvcm1hNWpcrpbGjI79rwtYAz7dCuUVJo4gSPXfqA+ARyUS6PIHYipQ2h0KcbVZsbeAJAGea0OrZ
pMwp/CswXiB5MRfkx2lnz9v/4gFav1lUI6gVZe6E6zL2IPoo2c+Jhs7GraHmpb1fx4BCID5JAXpv
9P4SL2faIrg5XFs2wlX/hSu+3ScrWyE0u3NOh+WNGQ3tlAv5CoaQ65lrxLbFPItdJmsDqWfZhgW5
BKracxhFLrfL4YlkzocIjv/VbPPZSsquIleA97fqO44s6HNE0x4lnIdeoNeMf3cBDY6Q9lnfVXV9
nTZjsFzykj7vjw9B302E0vNpb1AL98eBrUWdR5fdKDb3feetYwWccVgUzY4Qu22508OllVBhlmrW
CdcqfL/mo/W1XiJKY6hnaoTc1H6I92Bw8aFNv+58HY3g+IwhHJiFUTem1smJN5LyqZlsv/Rz1D48
3Ybwbysy392AoKVwVei5F/80xzc51u6g1QulQi0BBLm+HDBToesA2bq2BWvAVg+XeIJSeCf9Y9qw
raVoET7VoknuU3B79ZCtoOSMOs0017OrngDDPl6RVccm4VrjJ4hYy/t5FZavYQglUBhkliujDaXl
kLKRgTGJpnTTagKkvWNGwdEcpFkudo1e9X6V6pnAUVX29Zx8laFqoeWmyVQ7kj7KsX5HwhYG2OF2
ENULqFP7yBvm09gPWdWZWVkyJ14+ZbOKY9RLzHwpYnlzLTtVNR7WCcGILkrmKuCLdgLKkGa4Dbmy
0r9raVaUIcnafaXK993WG1CF8eOa5cTuLQtNlwLuzL/GZtkGolUqrDPsHuiTICCc8jsBczEwR4Kg
wL4QZBaOAfqNaQxpYUsuQpMY5IRFtRvYiGfeVFistNen0BDUcPUV1u8Wl7JjgtQKfNFb/N17xIfN
TH5CatVnnLtS1TZG4WpFPFcpOxjwzQXPIBmEKaG8S4Am+Ck+NcQZoUS4CzFKUz5CSO9MMRqaotbp
8EH4Co66mRqVzHfmoO6FWNj4yICUPmxK1zXAupJ/piKtb8lmNbPqF1W/MwyU7tWw6Jj8pzyQTDRk
2c2pVZORnhhUynC0YkN4rZbdTxi7bVLB2sCwCMWI+UP/zpJckWUMS1nba1NLBYCY4PupzWMGe0/d
ugwhw8s2loWqP+fHfuNNH7t430EeFPTmXxyw+Z2PfAd/tjiKzooU5T3aUFPN2IVz7Cx+8GRfPKBS
6kz/MGp5z96pHKyK7IyQy3atdZVLEz3/DPtd9rVmONxK+QZKx4KrspCuj6vjxoqQpWcsOiZBx9+X
QKLUQWR9ic4qd3E/OU4UeqGd0AjCm14vLaFQIO30dzcFed2JJaFLg+lWgpl4ul8IZrsTIUasrVXi
Bi4sJM6Nqc1m8RuChnofcF74XmjdmAGv8osY3mB3744eJzb3Xh18uTSvXEzYgJuI+i/XoUTy41a7
tHqMR3Gp+iczpl+42NPczEH3w/crf5algYvF91bcuRYRc9uYIp+vmeHIkCI+mKoxnXCIk1jk4jCL
dlGjBPuVqvmmpKIdn9Bf1+NKrAx7+K2sBxk8dXR9KLX5L4ql7WZXkpD1aIWHHAJgNZIj1K3JzCoo
jNzo0yaw0gSozM4J3faeAmv7zgDhvUubjr1x44OTitlG/LyBO3z/oSnmmaqXnHBvwf/6TBtp15fS
5utSwJIo1hjGGQUTAoqmBLZARNIAo5XAGCx0j9UHkeDvEptn9Vv6TdCVpXJuBVn1xR0qPki4QQNv
Bv2PNX6ZSBSQfJSfl1TrZdo278tlryRkRDT+J5U45FmzA+amsGilP2GMFp/y2YNjde51V8ZHdrL3
6Rp0PTzk2NhSbnevCTyV/QkfbUSiiaha6x04Uc2AG4mn85TfPq0yuAGbw5qVbtnb/WyjnMHLpH/j
ZccPFldPt9scUdJxbmFsOaCard+h9X5Hyx+7OS7gVf8GZoohP0E4qKKOA9cpxbKvq45iYjSDhWu6
g8elAdQ6gAqhYjqzdsGPkSW4dHWMtrC6vOXlahE5HMABHKz/4YRywcqPAu4PytinX7yKR3Xc3ubS
h9XT6h3CpdqrYn35Cm02FuryWET+mrDQb9Z3o47u+NdjJv9qh+rg0mTbUMrFvv4Tmq65Rd+bX9Dx
PcqLHGIOaWKIGON390hKnDcEzAgZMQbGsLidUzuMqCCsqCzbU0u6v+6itwtvWpO6jNnbVI+j83sI
IOFHlblrDHP/uWGFEKwrhi6wEgivSkSP3tdXREd0hXQKwZTK1bmgkODjIMmoDaTvfDvb4MGG5yJq
Ec4fKPwihjo7n5DqThuxdU+KRWm7F6Hhkwe7McG7R5ELCXXuDR0LJB5a0/6Sq8TOHfICd2GPliVZ
fFPPnDPDeh7DRlOUWkHRFAdgzH9bVFuliHXCcHaD14XOTCPbyzcBvpMS+DnMzyvw+6It7uYN7+2i
JZG1ErX8BsRjpJABIG6FDJL+0jupBkcdasTPK4qic10z3V036JCYBSpqoo9DWhjHPzt7p1zb5S6n
a3jNCqK9PpZrgmdtonlbcTJ0/FaWlLklZPy8QtBBgyh27vx5BZGLfQF8RDXII/yAJVZQ43wW3ByD
qd3hkGuK7ya0c6v2Yqv7hUwf5t4T0nXp/IBbcR6aJyTjyQGO2JY4Oownh8E2Spi4bUt5hn8mdw6l
qReZYE6MWtuR5JsAGc0LfhuYD2ioPjDLV8pCymAablHoSKorlEwKrq5NZo3FhOcYNz9Jx5s4kPhs
shRJC5sLGB1G01xsKvW1ePGWHhAPQu7mTksjnG6YuuRpQsGGnWRR+fq6aaBLKnAqUvm/bR+LFKJb
kBPWyaE9gFIAu5ljzICWr5FcK2eDfv2Lmzut6ygbcsHGYEmr9J1MnStM8XDfBotQrEBfOI/dsh0P
6fYX5RPaPiMq9jffm4ixjvWlip0WvBThbrK3Cx2zYd0CCH63B/8sNINB3d9KehZkzuTDfvl3TPH6
PzXGOAXv0XwIgK+4r2WFaieNdHxHFD1nCqOpJXOuMOrzIBryPabFvo9ergTV6zTZdsaZtFci7oei
1WWqZhBzyrQqnH4pram034H9gzGOLE6ZSlYGm6bmWJqr/sjLa8Gi/XwQx9gTGLousd9a9XY9+2LM
icOD87/+oLFpe0JjVozlkRJVjpwf6KzFJH27OLv9hgMHGz+3L1h4YsV6xpT1Xffoi8t9qC7Pergy
At1+q1picHok/gvtTC8x+q2UNJnVcfvaA1xJgiFYR8F39Txzd6F5NL9VQ+x8P8rgJWs4qgY7oeqU
TREHHF4/mv6GEihQJwfjZl/7/eyfdnF85qHFyBI2ZPnaM1tRY91atnzybZ0cRR6DprmJ9t/5I5XQ
d2i1QazaRJdntzILt9be9Y6rmb8rbmTHJnpS++JjXag1kCvnC89yPraiylzSFxXfXvrhftaa2nA0
pZSl89ZzVBZrvCGP9wKprNNSEyrTYPtKaW523W3OZzDkN9WYxUjuk4kTN6ORFQ354qMh1uQoDWmx
dBuaBBSys3FmvV7xGRn1G9eJ+GBWjd6f//RVmDw8zBieTrVzBACAM0pz4TuqPIQULzqeGxk0qSMY
TjV4o106YcI01stYz9C3Wr0ABxkW3gXq9rB/MCTps/chBxAksbA/OhLmsN2UarpZ/vshYrflKEIw
g54u4bWtiICKnW+z3KU7FOuLrF3Ug6uzP0cF17N1YZUJZJdG3rsa7o3eLSNorZc+TIJoNWIc9z2b
7uI51qOy3xpKFtAAe3LEqceV1PYAD4sPmm6A4tC9NpOXpfYc9Y+ZB31sGAxPtlOncS1ECzSr3NcE
SNGI9f2pqVeUTH286SZDuoHDmswh+PvNWviTemyEIeBlQYYmljiT/QHiQZ2kc+Edop6eV3wPmeoe
WI/VtWr4/uAhpeOztzfiRNkNEG2K8VVMFzHZfz6d1P7a7+Q16oJAmB06E2Pctc6sZSrFs/8wcUHl
JxOMKne4zWQWXpgeB+mQtts2mXrwrszUG4bpzg/455t0uqRrqi3rc5vJlr8qXDL4id5RYG6+CrhU
c5zRvA9i4hmiIRGAJPPNOlcZs2l167gEdimnZVRt7/TVT/Lc2AshYlUFdsV64repWkaIILlolIMd
aXn42NHM7C0ztv9HQJ/fqTAAsACrjkVtYwLmtfhUDWBSqU096c9WQO+PI6QTrG01IjtscgRZqxej
GAw+Ebjl+Nwysq0m0SeSxoaaUEBCbX/W3V2+V6CaakTECi7R0/mpDTGDQDkq7lM6ZB4vUZ5AbLpH
jvZoLRBPOa3K5Dt2aJPWFyy6Zenv8B7z49qYwkZfUXbcCvdEu+K6BWRjBv5wKrzN0hregJOw77fD
cvF9S8knpkX4cRm8KMAmviliOsRK0Xk3Y+l/FhX34wYgTDt7xyXYE0pkHuVQznsao/O1BVKhtKS+
JlLaQeSf8uPqYm+qXXTNZ2jVv91JSeUBXI0HJxjNpiwCYO0AInTFSXna8FzmK+TTDfv85y6F7as8
++15D7JvnzU4B26KTlefI8/Ixgpf2tHaD++tR85CO/FJZWo1bP/LWr0S60r3SGLnJSRO4pbI0L/d
nxnqy6HmJpKi7zou3Z5+QPf/OVHuOmymWxhmyTL7cKGRmI+Sh+A72IfFQP8oSmblfG0Z8xDA/BU6
wqe3PoCX/oOsdfczbNRx9C9nLnkXCDZeXDG264JUw99PaLwDh9jS3MYTDF1/4LaGnH8HulnjkmMo
dRYkG5RrhAbY/tmbHwqNqO1IpwUwfprLQd1SdhFNcmOyd+P+hQ9/WM9OO4wDgtpuMZ2W26nf5DLH
gpTES1AaVbliuQY/20/7g59B08W5P6TnzwKTIzARUjZDDGBLxvC7vGCsa966OPaTWSN6HW38JYsy
+0v7RPOLhlWSMWQ60vXzmE/mwKZ7xYWIXbv+6b/yMtv9jS3I7C0dDMaXauHkzEwwWEF4gnWPPn2/
UVA32LmXVTXPJQJr+hQdGHqZ0eOC7KMLffb9KyFlaUd57lPLsULXA/fEhj8ZeqbxxWdzSrbD291W
C0RzoAPVp6TaXCp4Hsmu1P9BVofCtNapqNVxpeyjSebvYIPrXrIq8vY38zxJ5XOCtzdanFI58Z8z
/dWeqnvmWTD4UnFLOjI7d3rRG43oGPkvMTW0Ob83jKMx0X8HGzZnb4f3RUuO3CdU7Oe3nBAmEIGA
9pKejVWiwBYzVAZ5ovibPajyyioAQLjWPQhv2FjZwWB9QCncXgQR1miI2qTIEcIRogj+bfAL82S/
DmLbc/pdea0jpOLHnYCAmLnOLsyoqw6yXlOXt/bygU7cqjqSwDxFmFSDmxMOvE/zu7hILjrOK66k
ESwqfgsxpoCbJ4Lkl9orIKRa19hQNVyMO3JMD/oSHYAW/pnIzvvcggbG1/c/X3NCtLnnTX24wytH
XAYND/smoO94b4+QXUqqSLet7XqavEtVJQ2P1K+dgJtff/6cUbFExPXrSXs7ciICbPhD13OBypIc
fnqDtrINe+E1nq8qV99BMKcFdwVk9l+JsWjvojFad458HFiTePMhpqLKqzgQ9G12YsPTZ4Zd2jT0
yuYSf1HAI7jn5jonWvhlTeJMHH66LLLbho5UrwnmgHprwj1k+yaJ63WD6PIkswWDzoxKEQRuiYs7
RgJ3Aj2qxvu72L9ucUY4tRlI87V9uCjPq8HVR4bsP15CH7SX98Um8Wmq9KKPUxsp14ZIu3ODKa/M
o+og4SvD4wxZ/lRmXUpbgj6oEGJ+qKUWt/3SASFmbke/7DtgnnXjIYHOIrBIIAN2ULZDI6jBSyJy
ibx1ACTzJFMqa5aHK0oczCQ++0X/exECJeqV7mTEfoeLtFoQbx4MdcKBkOTOrMV/Ymt2xtgBvCep
sYacmdNibUk0WnYoKzfHXPdDXjHTWvYX98RHTWADofCF8d0iaDp21Ys83kwQ5I/7t1WogpX6zplt
XUxz+ojHR9T6ENEcySXntpq+bgU1Q8WWgMCCjYmyEEnwr0KKTYJMs2oR4gu8wLOOxrdrgmDzl2d/
GhSFHuyqnzC9KMJHzT380o3GZRc+utQRlX67FXbIwT3wXeQQ/1TMxoAkL3Dm/3y0SmeahMr+qwfu
8aoaiZSciWEv/eJSRgcro7DduBaVLVPK5X7lttK0kSJYS40V+Ck1hLPndQ7LIsVd3GOBlWMylpF/
2Ipcx6/KJV6x61BUbV2jvfvod9qc+ORGUR7teMQe5oaU5Dzstl/F7DbEoV8BwGfCwCMz6Gix38lT
Igk171nZGGiGAZq6cUtGGkOWXSwpJHnWkMn10Il6oWUx9t204KNBfqVS802qYloYUze1C06YiMSQ
2pWkE/KPpQ0vuqmL1pWFeuDiACbJ9EBEes8zMtw/k8lCMVVt/z/QqXWYaibkHy4kQaATRFsRqcEC
nULvqC4oyP8GUFL35Q/WAKvFS40x++0UF8WZaRADkKTtgU3QyuzIi67Ed/mkppX+zWHnBuPtEzxA
OrabX78E8pA5a3rCyDHOHPB/GhDO9TEU4ERvs14gis6diXOg0BQNFOHQSLAPibCxaolP1GmQ0P7v
xABfiDswKv4L0yaBFZa055bZjoVTSV+4yEt148FtnKxsx9n6hYyqOxoWcb+SW4yjDWg6bLtmbmvJ
45VCBGbcOci0rBiDGidosbmwYp4oB9rv+5UM+QtvcsXvzPYWnzPT4EluhMJ+66D6MqIgohyhkCJt
ZVbCoXedhJlFl9s36bhGqCCVM0PkD4Yub8zeZp3o9UMBG0DOOkTh37pyU0AM1cl19WTtYi2vEscd
uUaoGI41MHGhfPMpkZAcKl2PHFQjOKwj/nOep0VwucGBLWKPgD52jflTsJ/MckMbQM6JngFjoifa
pkiOvrcelpgtG8vOaBxQhhq1BVDMHvo6lOJTpkn+I/2U6SnfdPrtgn22aFbPMUf4fggrzWAt7EL3
ldVyhY+QeAMs+tRQyxAyKe+GGLzV9WXgRIIbVsDFxqObWUYLx4/vXCPUGMioxWD1tEpFIk8Ws4ZI
Iu1CcTxCMy1ZqV5h8Xoe/zLk2wPCiTFrwey92qet/BfqeZT343cdOLVbrxAlkyY7F3pTxLob6KPB
OtvtS8+braJGWzjhHKa1ynNQ9tRDfIXR+O5upPDPUl8xNYK4LH9w7JAyjIzKqLyRFp04qp+Xhgmt
YGmdD0WQfu+lRw4/zz1//cto7YARSSIeuksIjFVZzGFWT9jC6J6CwbAddhCxpA+tignEzWfhEZb1
+UUjMzUZhiG5sRQ6sR9WxgnyZOyZjYPEnuFy5aMYkw+ltKWmowkUP8wI/p5WrBkBPrhgw5VkBO3m
Wh5GaR/wZKTP9Cya9rcR9U0yLyNaXVeHe1oK3SiABKbVJIif/QpLJUSrcxeaDKL3mW1DGkt6TkBN
C/Cnn533pBbhSRoEDxAu9JMXkyrxz3y1aYR/cwz6jZ4OKFuitl9IlyuYvr/gI31RXLnKQ+7GJxR4
P6aB84rDjBtHDz72EYj57SlCOf8tCV6S4cG64ZbS5YiBc95hmuwOTqi527KHHqMN6peG1nH7iSh/
SGpfWzHbd5PLQ+6nuLIizxHl1pk35HAuxxNHsiKo7j9fBgDq1+XMxqAxP4KHsml8aLLrOPxDdE+V
WEqNMNUyUWtVcdn6+lRnFINdE+suelb/O7ObPCCskG9QfFPBPKS81gsW4+g5POs+euolInpgcXwQ
p7x80j7UyhYTkSS3HRy2YAbhJSrwaGNC7SBnF+HKEZMbhA3efdvJH/yZHr69sQefYIgMcTJ5lEIB
ggJNhN1FnJF2q/b4Fg+GWCJip7Si3vjD37N3TfDLzkS90+87AbxDehfSPx5hFN/QOZq1gcgB2eYO
O6psIWU+U6glvQ7D9il/VHeYo6+tv3eqXJN9PIj38lYdB0ZtHbDO7KGrGm9YYV2acVpOHrtbbfSi
O1k+D6A5PIYEGSjGkVLBpSRP2MdRO4lX7Q/x4qqSr0neXWAuejLY05pAidk1CMJX4X3+zR7XmLXq
SCF0xgx9HN8djd4jCR7S+/+XN2qdVJld7FaOD3tMJniSiphAd4np0/dYiDkrx7U1g62HyTlf8pz2
ScQZdPL6IiBxgj7Zb5nWZMTyx3DZvM3GdUdnaG7QYdhEYa5bcLB6K9CYZ15BjcpfTbay8avfhqY+
qKbgza5vAEzEJhkL6hJU1vlHRvWMIxjnpqIaZKBJuxBYPYzOhBbLT0C6SbnTB/rnZJQ/KzUC6tKl
Gae7z4hV/URRMl1Zo7DRtnM2tB94Cet4yNvTm1P96S8cEHTIZr7Vu58qsvsadlmqk7TclM0SzmC1
JjG5tX67yWtizSYFuY32nyKxZkjNXvMFIYaBIARoujZDv52WPdnjtRfJJL3MINkUf0Ik4H1t3d4c
8CaA44f6Ir79tSxnlRoGNn4wCfusRgSjU8jTtHn7Qo0Yidz1PmWats2qcx7GXC/rpj2cmJ0TFSxs
B+KSLZmzd0nSPUpHJu35Gmx+2V/S4f/LF5d1+wrLy198vsbp11Ih+QvXrIozYwIq4J02xvV042VH
nDiuUTPcDj7MRYXhvWaP52YQfliRYZ3JA0lcbzcEf3Wu7blCbxbRTjvxLDL+tp2aq8TpfxjLVYio
A/+3S2A0w4BpNHAh8MxRXG5WVSSYu1T+6oHF888TnYiBZ23KZWGzVeNIH6J2jsBPhWZ+HypFqarJ
6QBgCM3E+BONpC9OXAtV8QCGQxHSHzUUUOHH+RVxDjCPa5XoNGyJ1MWf64/vUkd8TOotZGa/ds6M
e7UyQof7kQotExR0eNQOREpC1CQY4kOmONmMFWaJw2fh+7ZaJyE2HYsvqPLNs4dNI2uRq7HmM0Iv
Lh7T0+FrlWa8St3mmIs2jduZofkqGeipef9FZHSqJX7679Tg8NXacAqpaUzMXtWhRoLrYgPAxbh6
B3AJdOvftuhXy+h2iiyDDGtwbvW+BFXPnv0PY+F2Ruvo0uLb7AKeGVIGl05MfA5M0kLdeIeI/uGK
wMarWavPrbxGAEF5s05AI382eLU11hwr+tK/ZgNF52t3UPibwcjUfXVIccfIh12PrcocPzU9a5jw
iCT37rHf9/84LaZ5W3/IKZhRFV16rFVJRGoqUHdC3WUAkjHwUzeBd3oqihlvN58ni9RYpzVaiotv
poZpa2U98LNzrK+NTMIKcuPmJ7VA7zs0WeV7yAAMgbhiATZ2HtgnJ7Ea0nvjrSDBYeONMc67t1nU
VH/hfJo+fFmbBjN9wE8z/ZSmAxuqgJ6FjEoBtnZ/GUHNi2GPZvo/dOdIxLBD0vTepBtm/M4amhCj
5y0SI8SJD/pKZFu0Lhzn7b6S4QnbkcBaibsr+BigiauU1ogcMGwTo31MP4nYfGc/KCf6vfAgUDNS
srg9nGDMzmqXNJ4nLmfrVuIz9Q5vaU4Scka0qOIQUlpURUbS03zM6WwCafbp1itpMdWc3q5o7eNE
jqo6wK7VX+OM6mWIMNrXJYqJxeKCbrImrpC4DqCXWm/iHA8VHhIar7rJAwyaTYkjx6RwBWFNaFOV
j7E6UxbqJIr6FD169V4OOR0PXZCc7WSkzDCyZAuH8N+WVMbFVYeplCKU0a86r6wFtYeId4b4TA06
1OTj9CkSy+a3aEnhZWjFqi8frR1AEsIKPI994TWtyqx63/XyF9Pfglmp0CsfpX7PKc6rVZKDArDG
5Rpw5kzvACeVHYfw6+/P1h0uns7f48icG4+Gy9WA58j3uPZc9Qald68ykpU+1P9MrCWrYrjTckmW
vjflnda7gixuPFkj0OoRjTOAq6H7Xeo9HO2YBc9nP2fwuKuZ8hjO0FFJIK9jMIh5sB6ZTKeLEjjH
eNJKMi9Fis7mzc0n77HItU1Ox3Tjr2cMHEPZsMGnamk5ROfxp6cTvFT/y2vy5j4bdwTjIp20vQGx
IknSZ4CCVh05hZ7FOXdFa3mmaWp9FsmmFWi1c0+Q5C8/21hItf8/p8l6kRFHjaGNxhU8Q9h0nxl9
Rm7M9wCH9NTbHWjvmu44hvNBpvkDflhY0ZxIoABZltvNkvWGdtQM2e9J8Ua9TGfA6HhzV5eHqRc7
CDyMV+eQTJu72m8iqb9EHJWWQ8tr0wYJG/cfaJa45pOZPy/pZgm3olzr5/2YrLlaa4HVF6rUvLTA
q9QJ3Ugjct7HYX8/wsr18czF4AZ2FBpABQtZvTh+muV96qDEO+2dgznZSIqaEx0y6fFbXF1Mxpzq
mBsxNFYeNGBHGd5xABJ/dtfjUY7JN/0WP0j71IfuKvbC9k/9qvJAfowYPgXHwAJ+wgggO+MiP2/r
p7/uKvUcCN2ALTX16HPDt5/WZxzh6QYtDZqKi5/gPqfx7qd/gCiabPnYEVsj97yVFeo1DUN22aw+
Vut3VdepXYvAZm/7KlnyJIxthJySwI1mcXEKBHh6OYUkFOJZBlMhYybjcABbrJt3TMaCG/tLGwwA
cdHpDAW4PY1wzkzIofTiHTeLsmuA6Et/Nkq0Ln25wAHIIET6m5FED1mhARdGPi9Ia+rDRxDpaE9G
eYWNX0FWtAa05hi1xRh8vM4YSqKtnTEyCBD4SM3JU0hsk7smSZ9uD20k/8SEaGcXAu8xr1oc0+RH
PkPUL3Bgs/hmKJdGs9YWiRAOCyMb1pYWPwfuJQLuosNiKPAEYTygXgrYrwnuX3SwVeB4ZcfwwApZ
X4Wi8q0o+vV9YFKGqiecbm242rRTER7xbfka/I1kV3AP6dzpBxFecnaoHOuKOpHrgYwylkyR5n8s
HjJ8YM0avaNeA18mHU2T/gFt+d0dFP+vRYZVk6jUDw9kHmyPteQh19HLirsJLkg+N9s/ts2uKzfj
B21QoUa0rQSNVgiGwEKA9i9JE+D1sHHyYe+FLqCD/1iJw2qlYD3uagJ40ahXTdq4f4CRlTtzf3nM
Fm25HvPy61CxL+uXgpKQEQu9yK5xg/JUvxOGwM2mlPOoybnbtqN0JE2pWVBy0VXUF6LPmlUImhKO
IushrHIai8eDwSlfariLBuM4LOvnqAhhec4/CqE/8c6S5L28DXtcyW1kr9WXmmaCF4LZli4dVEpd
fM74FppAexMIQataWj0uSRDnR9Je08uhO1DSXTpbsdGi7tC8kEXSlF6axMSBz34aBhWNj3mg0reh
IhjZYCQ4Dwq5skaexciTAA6jg9AZXuJDv1NVkFfTHkiDc/AulcZSZe7KpHPDCdR0ZIBdqNRJQ/Vp
xxexSdFr2VHAbfB6erEt7PHTmCOrPLJSCII9Qh8dJdwn5LpIneI69VXHsADB0tOqVWrGMtGF1u1i
jTyJm1JWve8uOZls570/uCPEpg08RMfpBxNLj1MjHhjF/j0ulbwQ/Bw4jyq8U7f+3HqLyNzie07a
Gomqt8mo2ORuS6lNG4pUCNplQW8QKlRTdj1YGUticaxjzjsTaks3StZmO+IMYbBbhoh41c0htQ4h
jEvlDSsxH2vdfIY9uQwCR+iqh6duj777GHIYDkZgQ2egaFRZ18X7e9LoH4VKzfZbWCrASoM7vcG6
A5N3B/dGphP+TFI/u3e7EwRu7M4koBVef6zvrNNOcfqX4TEoDKiG0yIyMgUK/NhR7OzDg1SAow4m
8yjAEoutW9hIuDPIH6aq57g/tP1HbI5pDNErDOv8v/SHn971mR5y1hDxaEVzk5uKALlo4h8q52UB
tzBCJbfxiPuWdgqMky5w4NubIcULQw9qryK7E7bj7p8Gpn9jQc+kn8kQn21bM1gE5q+B/V7JRRe6
GFhcxH2H8EIfp24wN2UN9yX0QmbsEjD/jKhZIfhijrWKu7h3ZB602DTBcbDy0KaGD7fyd/+oBbBP
Uwi2tfmH/NlW68eStfNPGs0RzgqHPd7+IugdUCJrH4d/Wrt5zEjx5MclbMCzjERSQCbZ1no7hDhh
EYirMWRrlMmktckA9p8MXQnzQSUK10UhQ365TyetVdcT79557ZfZek/aKwOHgWaLaA03AYg2dLy0
DYoYY6KyKlcB+cV/USFAGgCLhJ2pNa+08SN52kqrvhl5ff0/GdFy6ejBVT/Gf6RW99/6qTOZ35ni
ZP0iQK8u1sZJBBjsDXGwL64E5f+QHBPIjSOs3etwQIHTyv3xZkEECv2ebTo0fo92lIwavA+M2pEp
TJJND3xNBzkzVB3IbLiTQYLWSCgMX1WRSfU0msaRh5Z0QRiwqDE7SgLEk6+Va6rhOGCSKcvfTimz
F35Mo/1ZGu30sYXaaUs5JUcHnnkB9EUqVA9OwAJ5jcIemFhHx3yDgOQpyuzKnG9HZUVI95PcISmn
H7ZkGqXVFn/jG+OugNpxrSAWt5QlOS14QWhlHQMyYUDgxxB1jvqdwyE4Hl/Nr7Opo/DcldOw4grO
iL3ZMQpGm1AFOVXwyO1YhiUis9c3R/1DYUKavtDAnsYvyM5DRhGmw0G6riPdQNxA5v2R2w2MGhF5
JVRMqjcjLtyM17ZKmeEPR+oNIrnPqq6fikC21+506jBGunavE6ytp2U2FyxE2+1DAF928znIjGlg
zLbrK41oPNYw1wftEX27egV7HjZANppSrgly9x/M2/tiMghogWwaq2jzGnuU434FxAn7oEGTZtrV
Lh69MtAygaSlfWtO9QNBCooDeA3kAY3+BL97C9xQfB+O/Ne8AHJMnYQvZQqT0xCPmTvhaGLMF2oR
Q5DOh4EI/TWVLyMtHfbDk/PGX6fddKxShe0kUV7stDNqYE2yyO1KkpjKU177f8qGvkxLKEnTtXak
Xt0fvP6v1zMJxhY/O3BYWA4blckVL4qJL9shtQviK93EqvGfLangtrMMUzdtTgTvbqA50IIWfeMJ
E3u5LsUWhLJz+Es2+T01902KSZdU1IW+fVHLx9brBNg3+vEjJZFXb40JsA6gGOq0mNEX1gV4EFBc
9yQi+l8GqKrM+9kEHlfbyszUJSA9CPGc4AqesVogDKa91iduVXSBdOc2huEmQe3KaKnWLnHcoDoG
KvUSuzNtjGXsTt/UMI0MusGYqwKvJerAHq9W/psfEpsBYRRzG2aDoYhpbir8kzphvXV6CCVtV02h
mVv6di2Z6WWKfZzvY8NTU32pdbhhxdX2q9e6L4C1HVGcWmUm4+W/CMYqB0mtjPtrJ4SCKPOwj9Tw
lt1XqndzRRDVIAPLxcLzkP/qYmN3hjzU3SZ3wJz52FrX3cIcuwpcpTX7CFls3F9+UR5RCX2hF0zS
2N7Fs1CdPyhS4N7x+DhpNL5WlwKjfBypAisDBcRZBcVYxZZTgcb0Ci/n5ihKQuMI6ILbZUasYQgE
QUB4EHpqM516Atx0AgiMB2v6UbwF/CNHBl2foRSOpms+gL1AsyvoHN80QWQRIGKvpOJyU22gSrpF
rbd2pW5tzg/Qovh3QaS8675vn/uhRipLpzoOJ+0nzNV7+kfw5kWuLscwBhyonILc6kS70ROrrT+f
SJ4+CL58OCgcf/dlbbrxsuTawTbnxKvrLW1E6ev+Qre7gradQHd0+AQSoRSpkvcbwU8cxeFbP/MK
gHZNRHjD6r41kl0iN0U4/HO1ZlF8tfnJ4zKaE6EwJLaDjhzUcehVaW33N1EZc3Km2eRJWCeZnndC
stqT+HZHlsC08eMGP/HSYak6cMPSihG4yD8yvzT29Bh9HPvG957l5WOD0jcMQqm0JJixX6UWaOtX
s/krZMbAnq1pD/R8G+GVpTA8tuQZrPNr6cWufRM8PyTcPFsH3kqzk6qrbcgNKTs+nr0R3xriCHmD
qLA2JCCIy/slJ5N1uSa74Ovs8ml5dzY65GYp+Db3gcpalmQTJ5ecf0xVxkaZUnB85vFvK++gehfa
Q9wfGiopzREPuW0TyzC+X2C3yCsWHTtY2CkagPYtzF9n8WxBQnqAz7wJ+LEo/S6XZZnT7lHViBar
THyNrZk4kKzJtr7p2M/yTFcnfnJdod3TX9HFkhhQ5YGw5O9HBeLe9LMF2ASDQ2kuh4imUP4AQ2s5
k3dc9ZN4J5iT0dsli7N2rlmxLCABneHO6hBAMLNPuv15YfYudJv0ah3JwfPMELoAcJ4tJzwOEU9B
0pFlLpStfmc/sVygpjpshd4y25XttVOBAOYzOkryN4hCfKc5NSf/W6Wnhl8piXrGfX37TN5lfyPf
AZiQ2jyhAuuvunx/EYXa0JHH4VoxdthU6juMsFGk05ZEXOTW63LjIE74dm/jbXTjd1A+d9swtKFA
WfjiJQHefgpz8MIbjgNyG6xHHxw9IYCs+WsaBnTmKn4J6y2fcAXLxGwGaznA794Scpsln48u9LTC
PAtpON5jUc7nmbIc1SU/yxf+/oHRfeyzwWYAuiKtRRrLU9sk0myDr+3B6YliXQK3Dao+CQg6UYh9
/bvQH4knn2H2aHRroAWlH5SrBBM6NIKNA4mrcnsrfOmqqaZyn/xelSCAS5QAjPFk5UyPeCx1U9VU
wdWEIB5B2aVNpu+owPXGF5QMuPzEqmIr6u4YTi/bbN8VH1fb20kT/5nupAzym74FlUH67CqGo2og
qDWxjXG9cDq77IooCkgQu0EtlRt5HGN8fjS3gJZFl6l7SPmG7tUgKasD0qM8ZqnI8ItD5BW08c39
YbEpFl3Bxz2BgQmdjc0WrDgeDl2pVS+9w+4yWkyUmDv5Vs52TsZdpg9l+V5QnY/cyMPB+X2dlWV3
uigbrwB+AcOI+0yDb29wP+DYujyqRICpYx/bb7Hx2d6zlda0scW+qkgwvvFxQanzuGXX9NppXT+K
mERSFQAs6elFQtcS02bdujPR6WSxx3VeQ+W8rB1yl/tYtQZQTMXfoYihatdGschYluTAxVLDeorf
YdzreYs7qwNlcaMeoI92mApDqzjCPM0kVKxET0iPlGyqTu3oUBeeIT6fis/zQHT/Gwo8ZKCMsk2Z
jX1H3pDew9LcFLIUOs3blA5hvjJpsSf2L6GeORkizNVyvdxDZNzGqKKgzBe88HWGf+KOjYrdy47y
TGVYRZMcohju7uIt4hQ6sJTepM9ZWY6KhNZSpKq4Oss6nzGyMYKKpoGeggzF51VWDbUnarUSL/tE
zNxdtbfL/3Ae5TWCxaEElTEuUBBqq4aN+3uU2iS/H/LPSxCHoRAvpFuPx4YE1u5TOvbPiu+k8R5d
ZYK7TcXYdmK+DFuFpbjdpyRdQVGt9oaLwWVCr41nrC4+7GsrOYI4r7DGk9WxsdywuOyuCQak/fga
gcVJ9qC+IYdeUpOZ3ytKYe91axgfyXmyFJzWG2CAYyEOseNkaUN46ebbQmuqyiRxEI9xtKSdhNyA
AjHXtrkIv4TYqjxiUzJYLmqe7j8gmAB5HPFg5qgGrbwy6vZjHRz12y8jcxtl/k9+PVlVmXEcCWKf
Bhc+BZR9skr64fTZgroFyDHJxyH5j7OVZJgy7RXBsQFkoZ5Hdr2l/E9I+zxX9nXCZekM/7lxuNEb
eQZmmwW/AUEjAOmE7Zmc1uuxnBkrKT5C5Ui4dqw/FxanAoZYXVukcD1HK7/6eAKxXTPtj3YBbJgc
Diu+Vxqq2/ufX9UGRlPWEB65BZRn9lm1+udd0G1O3IcdRcQW8sUhy6hPMRi+/WRXYxhgrkahq0LJ
UuzRqa85txYGi/1ry3TFvK0W63DvWEJz90zP/RlA3C46WwtN7P+Kw/1n0BMq/hDY98UNSa3hFH2k
26PyzEV4l+aAVPk5upgyxesKWphpKomo1P7nBpbX/5zjhTWe/RFUubt0RrEwP3OKCQ2IA79HgCyP
m3LGRzi3CLPFdY99RgxhlsRyfMoLuszbaQXkUFXYaX+bji1xks/9a3meiGGumJVKvsqxjCC2e9nG
BmW5g9+4IHs4+ys9lKKVanAMHPI/wg/UUn+OAkZvKY+LYkcgGfvAKZRS5VEGTLAAAISwzPqNg4NX
ZUfM6rDoh8bUdCiAvgJMIc8RKGI/W400QgKfy8LVnER+Zhvc5YPYlmbfFtob1O861LM2OssA9Nj1
WMGB4HTVQYzlxiH7AbYFZWTw8WqRrmGxWrF8V06p/xeZlnF4DDSkWTJY7zEqFWI6bfbK/TEhaxkZ
ks+cJcL0774kW0dKDY2KP0CWDyNHgBWWOQ3GB52ygPOWf6H2M9ag5+98vDHdsCY/g0w3G9o2bzfj
zLvp2YzWpiOr6cya7tui6/tk1ZypU7CJqvqED0t8IMKJ79WLYF/Zm8fp818q4L/vOtoSA7QF+sh6
SSDIT87lnV8MLVp3EMcD8MGPI9Sx47Ve3UsAKQyxswjPF2YI6+3177eIucvEX/Y0rLSZ3qzKJwCF
Gq920iRDJ2WbsOuaXK3vtrkm0A3/nmF5P5uDD8FjvZps6QgFnXxLSENjUjx6dlW5wi0GVFJrOXnc
eq1xznKsrdmYI26RWdxb1Hj0d1KERaU6b2wO4FRcFEjAn/PpIEzh+1osa8ES56W7wLR/qyM8WysU
PEmCzfbb4+jS0DujCI82u/EmvAA+LYg5GHwrJIq7yO3Ypk6M7+2RYK2O5V0Fn+F2XBHbpCk0aOwd
LnkoVrYacaUcdex6hmG4S9jKLeiz6e91Phiy1eJbbgS/HYtiryTGsBF7d4pQUU97EnSoRlyvOjiF
XwwsY0DGb4MmnfVsiLzAOsOKNevfkIUk9PTSonuqihedI3q72W0OUt3746fPqqUIGzDCQ2NiaFmF
x1hpW0jOncgc9CvaW9SzPjslPHTIOugA+X/g5fVe8UFWVxULgnqKsT/xMfEkT9AQ3ceZMy81R36a
yso1CHaeWyw4a+bUdNpcrr9wVobUsyopcn2nXmysv/FkZBg8hdG7moEPn9AxnsLT3doJRWxcQb1s
KWhx+Ev1Bjq00JjNrjsDLuRDsbpCYjicCRuS2ySCU4d+8bpyZr9Ka/BVbqtSLmrhQHEE0i5XyI7M
GNmMxM7y3/EK1QlxdBWamF9BNxPc7Y+osBLvQHImjASxQNiruc27u7ibKDFFdywVCeajJSD2BtHs
+KQ/kBldyRLgsnKOkuxyQtvh8gB3tZaSu6BnUFdL5t6wJG3ymnWi0rwlV3Wfs4Fb7k+zyxFxhrhJ
N0uMRx93oFFPfgT5/x26e8zaQVUkaBAZ1o+mqFNpE1yf29I5Mkrlx72Hhq3Kx9UV+UM+gAS72mHq
D2YkWg14S9bk0rchmdxQQq2NTNea8lMOOPI+R3Eo2g/ACRq7qaYUc0tigYDReky4UjEcDXKNxBvo
K/EEJ4dY05c2Ahxzq2vBPbV7a7HgwfQ8y4IYAGIEg386yBSpaFePl5r3Q+GjReYbDDFAvD15w09W
iXghRB6lWWzf3i05+R97SCflasLzWQv+ZkF8g0O9hN5b/dmDzgifyMNhCnlmpAdSL34uBrhLslc6
CuaL4qtX6/GTfGu6D3a1suA1sO+TXh/GzS1pORedmMxHlW++h3widZZT6Xi/4E31LfJPwf5Tw0DH
mwbrb0k6FjcsKLYQGkPfcJOxCtBI8L1d3p2PqBPAk8pkiktT/DBWaJUGxRfM/NtW47J7QAmimxRp
L2eMBsBk8rOP+ViyM7bZCTwLak9kiVLLyM/n8L808jYInGRxLaE7DW9FR9oQUmiLA+WtpDYlfYAX
bufldhkVrLtPoxll137BmjIzwHtUVbzgC3ma0/6Y3BgCHCUazTwWxfBzBvZTZ/oCXJHNKLUHyZUT
q58kl8ceSvcArbhs73B2GvlWSwPVrtMBM8VdLxvF6jeMHLiE1NEPGd81waF4/e3kvS7gJurs9YQP
1a1/QFK2pWhe9D0i5mlQP+BhMj7Q1k/T1/0L1NfrUHTT9J4gOWu78TBc14TC7whroLc6YeEpyxMU
wDVyM9r3SCaWr0SR287GwfljeP0CbvlUdxzlKfsX0QXYFUciXL6OXxLJv5jl8SqrllSsRxXbtYb8
DUIVhCJfEbfrcRj8+jt5jENpuZ6uiV2p6Zi3OpkELVuI2q2e0w/OLjaXCz8/ywt1Sj2XmfZR6lXK
laGqH2Hcr0hUTPAUXDeiRRznsdgshDQeK6A6uOpwYu4Z9KvN5ITzUW3jRmuDlQYiABwTAQw3zDNB
ZwgF0k7IFpqnuWId7nBvDhN+iaZtUAC+knHdXwiiKef3SXhKqYFG59r7gw6w+siwiTqbFngof+Mu
HoEC/28XgdNnXtVdceYCLRM5cojElSHeQkYJ7DytvjpOovMG+lYx1aPWoadqfw122TpTNrgLtzuW
O/QYVZTDtXnUmcuj4607TWt7HAFqNM+9gZ2eXbardpuU8D+vq0xgJYdSJBWqoJrU4sfDhLEWhgbl
AGoWuWBUKRlirDaLL/NOUVoAi9tUi/iDLICbn7CoY8w9TQtyFVReIyrMBDBL77Rxbv4ffKFFFV0U
0S+RlKLTAjWWIJ3MLMHfoBtQZ9q89nzQYSM3iZ03N+6whubdHPqENjE0p+RvpeV68Q4xzv9WebeY
BDjVmDbnGvL6F/faDdl6rSiiHgPO1HrGFntsO2/5A64KHo29yVMN/dK+H3VZYtjwx4fmks2aUXAG
9OCnbE0O9TvU4NDGTWJiMcTKQTuNnia6Z0dFzXgWrJVkATkvdQjyuk37J62ANgUrx40ehJTsJXt/
C4GIPXf+/c7/BF0mD6Q/AfYXo/sSVQyEqLpbhGOVQYKb5I0MZE2JYU5IKB4Vkpgn19ACbKqesJg2
EZwESLfvB1Bqh+PE+DMXNPyC3tx8rJO8MNdwH+JRDcH9pJPNMjzX3yJiizsoKrrfuLLrBEPZ/tDX
Rqk8hV4mJS4tsPOYL1fKcm7cVyaGWriNXc4pKyAO1yl0LsRqoAEbhdJbeR1/6dXAm1vA/Vcts1jk
nhMGgVH5dGzlHbKw1Zprsa1kxYlD8AK3zvRSntbU01YYD+oNzSsLrPk9DQcfWU+EZBZWka2onfQI
xcN6i8gEQzoTTKwJVjvxSrjcBYWFkGWLWI7ywg/pbEzc0c9/CnnOZRIRlSm8LjsN1ujdv6ZxdWKe
V7KRqn00o2nMuuTLji6lNAeUbrAX5ZRojN6XOAh6JkbbkvLQWpohc+vEgGaLmt20i/1JNzFWRnrL
6H8nTrdJ2fakvbYvl2j0+2f8j0qIoErC+CQuLXvtGGgTJDLRlIDVwKVbtJkP7ZOuGLtxsqnRMJ1T
+Xvs6y4f/RREb8y3s1xmTDLx7aFUJlXGsUHkOu2DxPRxAcyhI6VX1ImqEKu+4EFlecjK+qeoY1tU
fzZuUimBYbm1lpoChfSHkkwdKUrIPLoueUlXWtvySWGrYe7dzMJvGJyumNGWo3EbieErro2RgQDs
em7O60p26Vbkvpiozx6q5ZpoErrbb68hF8A+4VscsFKx2B2KeZU/keCEzn8DUChjCt2cd8nQqPy0
YsxI9hBifqmVTmp3A7j1o0QDYcxi/QOLYus0hdWRGk31/YJZi8KHl6i88Xv1plDVMvAw5OJPiK29
yln+QEWEhV3Wg8yczjCitW63DmJfGe4+MzHSDBHnudiLMwuLEn6qpx38ceSMUCMenMOIEhDkcsAB
UWMFOTktUnBEJmVwOaSDbiNoHm2GjX0Msi38VMj9m7hGneDq1l0QRLC58p0BDjqSBE8DH/kci0RL
ssI6LftHeFfzXkayfxFaLpHKtbCtGveTGZV3EHktfNuKoiEGDoWs1/6dbeU4H86mx+n3rjlYQ7Dd
GNJjsnON28KE6Ao8gf62SUWOZSgeua+PbH8AEYwpGmnggQr+InPC6S7SpMBxOOkH6K0jwBWyjNup
RrDr9cswc9RajHKKoTnb96fbXXjunvBu5FVpv4TLR0ujzX6TO+9O7xSGYql5Pl9ZFkQNyB0tpM73
W6n8Horal9FDCXKq52vSjJx0g5gySjjnbCWEgJRN/HXXjEZFnR8ku5qzxaMzUGZ6Qth8MZPabVBF
vfYJksVGNxmsrw/oNCkxIcVi0uFr+c7b4cmu7ue8QPRko3SirDT5HKALUqap4Sc7EnaNoACelQad
pX+eHut/e144UjPF6MmgDFdPx0+m879gL4sKjcVi1hynCDPmCamoaOR0Ij40PXbfyGi0kBNN/ffc
D9Xz8ljkWvZS8YOKgNuPQMNeh5Vx0z8tK6efWOMd3h80q/2rEKG40vruYib1UpecqtwFrBhVSK/z
vmcZ1HBT8f21SCKKTH0mqlMn84SuLGE9kBRUfeZPeLRcoJJqca6KR0wMh8REzTno9Zgg50Gqwazs
7WKdJ/+YYTqcMigT9nGU+j2LQWgRchau7HzOvelgsSGJw1FXSpm7O9tsxjGlQSCEMv8G4WvKRsWe
HShtmPuXMWoR1084ZH5+dhWX6B+duTeNiAJvUz/GTLbDm5chXLSmOqp1M8CkJULQnTb82x4nRAmO
3lkRonvM8r1epLzv9Kwmy/WXoOCpuFGVsXWB51uCd/cDiopqhlQzVBS6rPHan8joWBGZ3r7BLo0N
reMxZpROh2J8guKz6mTO6yCEqlJ6XuVfT3aszusIF8O7YuelblSTF4NIcxDeUHrJaXz5m8wqFEjO
F7Pdn/9khK6AsNC7jldLRxfBeZNzOKsr2MxkFfGwLFCMps1PRqnDMqXu4SPNj/tK3bAhSB4K5cAa
QpwI0XBnHrXZkqI4khMZTGQIJ0cQ0l7WmXoGg1Eu3e2GAlrJ0Y2tXt82qjFOnQw1ORxYUgS0PGIv
gdrhFEqglbXIxnSeeCaSUaTuJ6wRji6jrNtofya0uZskyWWOjT7nR+UUswegI4z2rtklNP27UUa9
9WsLu0euERIfFHJ26yfOzV5P3LOwL/HBomjzzIZ6mXTJJOPuBuTNQzF6HRcXM1rYG4fKi2L8BQe+
H1X5pU8nv4Upxa3Kr9jrNQdp668bhGHSgdM6JfN3QJDiuS9f/Egd9q9tIBvnznuvbMQVWHN2NTkZ
SBy1WhNID8ZuKJqcwIkPg/n8YTB+O82+lTAbANEAaffXXEKR/4Dxwcl4zYFbATDLW9PVQhY9l8X2
hcy3aIsDOkx/o5TKHhO90Yagdu4MOvuF30B4E/mo2939QI7p0PoNeDKwEoqLP9aVikX7y5mfWTTr
kHu418nf6iejc0xbhHl9D+AvwbLdXLjDs5T5A9MjljrZfD202rOeSQo+EJS7nfe7ULVNW5scmG76
R490pbHgX43zdCYL64UBpSBLd5GqCD8xeoMNXB+qeTnQoPm4eYgrGFXc/YZzf+wUfpPfiyyPVjm2
xCSICcXKLPLBheEvm1boitu1fl8kH3wsl/Xv/3zHxCe/CczdTlh4mvc4ugpItqzWmjO5+tP0jMQ5
K84JKw5r/0EXGf7LiisdveOLTUBQopZIDihrNhE0FZXS1hhQKx5xjZ1mSb9O6SYp0VAAQZJ30sVy
llIMvBh7b91cLhY2AF/B6PHl+iKUKaBwmRLTz+XP2DYsaKiWSVLeHpE3o5+xPalN8WwSHbXMryXz
PA8iW3AZsQL7prVLvke9xewFgt0dpzfIgY02R6+Masm27okfQ1iFtJ1leB4IF/YW4smgBMG4YaX5
HdOPz5IeeWNTMLwNDDSpRagWcxPP+vmEKKh2lQGcaSJcN4SLLvAhG0igkFY/QWQjROmc+0+pG8Td
R9ySP/K84Os5tN5tUX0BeilsBpTaTlljisA8xP+Nu+Frl7ErAWeXxF6KaRTFZXgHLcx3h8XsjRaU
rknCtvbtDg1kUL5t3NUJp4wO5miFWaTBVIiEBCDDGRJizC9tEGQ//n5L0crVcu/cjaN6QZbtQ9OP
4TG7gmTnPWbHCtS9eZNDx86Yz70Dyt3b8bOj+3tMWYCOhBw/LXfAWL+3r1fhml1SO04+RVu+0Yf0
GO/VITGzmYGDA4FV24R33vl5ZbrvbMC/kVc4niz7sSDzgrLUWC1zVyBpBYfP19dyRlRa0WFwlqAj
FXXKHtwcdofi2vDOdC4Z97IBjvr5lnaAQBey+bc5VGd2f6q8h4u82dDSVHTbmSaYSK3XXZSdKOY+
J9/AKa6m51oqWezeSxRMmMjADdlRZNx5mQ1gIPilyJun/haBQql7D8TD/26C2KIqwZ0iABoH10Fz
wqdSNysnpHVvUPgLkgsRRyzrdCVWm6M7ANh8PWCr/BGIWbGp8syJ8IglmiYXj68eff+OLzbCE57S
8nHBKQh4PZRZjDUKTaurSVLyjHgbJ/iYCYuJSb/Df2gD5nqO4GPFH82jFsEsx1TjdjQByutTQUFx
tK30vByYg1ap4+WqgDlrNw5h/v6ZdnsLu7iTMuTm6uV8rQQnBzdK+XYE11jNz0bmPlTiUb91HJFW
lnAuiaio2Ea1dvSv/QZSt78SllXYsNoQv5I5Sw9cbNiAetWSIv+VZ5lqSN7leMNwrDS2MP4e8rmo
AZJyV//0ak10gon8KFKmzRiyh0no7lCEAWQIrQ4C/jqS27dcUNgfFeP2S6wJyjdMTGQoiieIOJ7T
snSrZbdBY56/tWafwPWZIuQVkFVLC9DRwNPRlgtTjEJutmFcnx6inEQE5iqB8CdJa3drfDlidKlE
KVb7ygUWvRqipnok7yIRLXJ2WbF+wu/iy7NumMLsK19SBn+caqMEBR4OFFjnT1W69F7S4lX7Jiom
cGMQbHqQ5QzLTTZrFAAnDWXEYI4YOJxhUJoj2JDv1K2QDPtrovo/BDfzoP2+BNnIMa2stOeF5a11
SdtWwUwrtb9/k2mvkYObHuQ2YLrNpLr2QmCvpM5IPBcgdlpSiqTPHETHCkcz4Om3hfrM3d5r35aL
ocI7qLXkb3eJnXP+hv6eTi8qmErTLMjsF6i8NhqKrxOBIRTjAO0+W5s+CfEWTpxoQf1S2isN/h+X
F09quvG/2vyMMRYFOJvht7PbrIeyIAizxO4TVbIlTpZeXvUF3C4VesoLejk8nIQNWz6G2J7Kbmrv
/roFJ6MSiLPxKYbMvXOQy4RAlRekzrfeIW10dD3wg+TzHoOVgvvTOtsjbqFX2CtFlRW9AOazADdK
y2HzDLvMGNCri7wd+TKZpiwU2LnEjIgfaXkWlhBqqEPsJ2YxsdnKUxH7B6mZCogUPrIk+fKV84KA
rro5DjZLlh8Nlk3G/PqM+CvIA4D75rXrJtBg+wVYowyxeMbVSbmV9uvN70Peq/jnDdI0I5L/0foA
ofo9frsI1Q2RvYRccbTbnAgHiiRRaygNbpW+wJa0px+67ebtYpvSnJqRfay8YNixpsGlc07rKU8g
T9XBGOV30ysGp8Q92DjXvhCL+A1o3bA2ygRVIDhG31lU58nMO/ktkpMeXM7NCkA2EtNEP5FZNGIu
Vsgkk8SkAX0EeoV70WmWYVRHNZe251iCN8YjvEIGrtCFCtmIzY3yADT3GHmQjlOnpibzBMqH0+bZ
j5lMEe8qyfq3Dl6NTTnQGM8XrpmvpAHv9E6KSWAV2wuaoLc/WBnx9DUy6mxiQUs/TXU6t2DDmZJJ
FVbhv8WAS8xgBdmhBTGILZDF2rzCGIU3hDFgjMdNn3uWQ4+hGj9ZugVd5xtKBdKcc6HDMn1tSRvM
iFQg72efdlKdTZXGSKlIE5KbHEPuTaJW+qzBPlhnBw2T5M6csI6UnnwM2i3HjFDa5pfWsDroavUG
Gm04lsLQ/dmmdW09jV4MOQshpvMjP5bXqNbhX6ABUTfoBa2hj42WBJp4vr20/84Am1Mdiul+VWsy
5FlncxihcywmTzGD2UcNeOZmgCJ4FPNIudo0h8ljL2K4It75x7k7qWY+sHRCuqlxRCJJd6pd/0oB
ZMLPPcn7HalSOfRJnQJG8sxvIJtyTIHp7lgC7FqWhzxrVoYvh2pIPPCFWKF8FYVzrmKG7Bwkvo2O
Haa2gXzcqvNtOgij+7bvXZrcfid+CVuX7zywMGJNnhZy35zsCtHEpBOu5PYercsu2DWGUiNFpSsg
yejn4wmQ54qz+WAaxkp+ZiNxWwOM6eq9HvRWe2m0SEnKQxe5Ebl6alueL7vtOw5gLI5ID8RFt0yI
DBczQz75xuATFGbH2F1ZJaWMNcX7ccCoXkYKPHC/hc9maeT6URBvVruDnDmDy1IxSRm9dQrnPkaw
4xsERfSEyzSxNFlUTGt0QbvbDsGPuBFrOT6vHTGSjfSsxBuXw6P7kHAgsjTHMYKDZ+9pte/7YpwG
2mCdqYpv2bJiduAzgLYbQlEmsFt/VyK0RT2t2fOFYrJMhF5eox375slkUVfHAaDUCFcNV8r9dQqu
b2N+D2+w8aaAOgUpLLqrFBpiVas3PhOq70DjTyA8tQWQQIuTcSEtn+QmV/brttNJmNw0qN0qG0xi
FVyBdtSRs0Kegn/2cLFSFK8sEnwexisWn388FXh3wMJC5+AicYvVZ5uJYCwrmaXVBmTzR+em8Inu
TYWfFfKUZ0FpQZz0sDTvF+VJb+uwzEQE/EQ/JfOPbGtJm9WxR5ME5MoIqWnm2gawn5l/k3XSvrMW
b9F6WfIqLMckb65eBDxMq0bjAAaA/GIrbIAT+54ObmjPk2cRnf1EwPbHLRaHCr6CCCs0Fnn7FRYi
8gkHcfz7JDC8NEBMtWOvUJdcr1UCXZKVLYwGUUiMKIvMZTaHha9+LJEQMkF39RXeNN/3omHCSIs8
mh5Nx3sHuUadZi2jHcjZSry04pYYRDkAy2NgdtU9Do8IipBcEygNsJkcUvKq0Sq7C0luYCv0fMFF
N1d+J5VTzVphCFfNdDX/6DLjMPXNvVlwDc+AGV9nKs0TTjsdaxwBcMe8GF78eXiuEQfx4rjsh4ph
LAbzuFKfmHvCVMzkrsxy/ezVlV/DmutUJTxv+7PZ/I81MhS5bl0nTVwZJVR10xMCLkFwftaqeJli
K6DFAfF3BOh2dIwHrHhwJQ/egLLB4O24DSxoChFKtugN6OriRQdgCST5yxSn6ih2WQDJl/cCKcqz
Yun7PxaZZDSixit5lakp34CT7AAcKkRYfbHzFHuBu6LosUnMJXrpGGrXgSe/zHkSdIVZYy42of+2
MA4XJcl/AsbRATH0QkUO8soAet/TDD6pmRnlIF79CXjPN60ih0HluoJYtX9rSFh8KgG36UMNxgmh
y1gkGGgI3nwY9OsbjEy/aC7afVXQpLUtXzykWOzgg1HD9xf5+I6CzjFwy7tmFxcLLbtr4mks28mA
ZRELNkotgZiI+DfbNEGePsbs50fARGxsfyr93DmVh4jZmxo1duVO8Cwwi4m4Gb4vgyNnbxIodaYk
5QUi/xL1ijbDR3tDWswn4QsYH05Ra06vT6qwCQsukieWCk7pHCW+VsXYwXi3k0JHujeITiMC5ICf
YofYtUnwcHvwMJTfnoZSNM5vW31q39sb9/jzPZccIGb63B0hhV0nKynT+LE8MGt/6nkdOcjLqZ/m
567TYqKnzgBfyDruHZ9jNZiacxZ01WtdydJSqbPJcBbAIWsbZ8zGNrIgMkODt5zZLFhgEYnqvcQG
PYaY6T7mTRBXr6L2/9osK5JRN+WA+8EdaktVkEg7Vp0n+4fJEDS0MfdP/7NF5vZUpqpVuk7ZihYL
12GB3BJA86/a65R5BogHoTTcy/CIvXe9NkPpEWa7uJ5rYcQtZR24grO8RDXzGcjqWt43Nv6+EJQR
uCnVZvEbcqBQJ5XZPMeTePJCMo+awTh5lojqRzwcWi59wQCCwpIUoJndwnRVuhXRA5qU3ktMGcDu
d+R1yINqWNhVZ15Ruc66umfa97RnlAn3Q1qOoDGB0udJ+df5/hRACDF39L3724Mncy/oLjzFxwe3
U8TjcM89AQTVtOduTn75pgGzWvFLnpufLsCo7ZUuDltPCokdnhXX3PsJGtYGuknx3lvgJ1fz8o1a
OqCjUlaz6sPGw6pa3d/FOrrNGJd1kbbdwELm4ieNODQW5ueVY45sSasV39pzELMan/hxcL+k6Bru
mst8xtq5n9YDwWK6xgmEBe/b7hPJsqKY1HsMa78qSDtSYjVNV7OLOAF8rBYVfRUCT+g6yS3W5cHv
sLCCnrKEyCrnVCxDRL37pUD4vKO1prAO6y8V5R6cSeVw+8qX9ZpHQ3F/uB3fg2CabnB7VbjBkK+O
5+ZJokjNI+efhOWlPubUjKHZkv/foLcgUL9T988DaVS//Ufzi/ZSkxkVDonZtxwwLdx9q1W6LndG
VLUCxFtEXXbMQW+BSuwH6R60rh7Hvrtc34sL6dsa8KQCHQY6q+zwPTooLnUNd/rQl/IlCxFw7CMm
oXeU/+K6FKZ7WuQwqq9tnzcHnZseFO0VBt4kZNxJah9VsImuhmTsNMzQo4mJrJZgkYHobJxO7std
qWRJj/XGO7RU3QFJJeJ7w28WHeSm1iTdW7/VVQjh4+sofJfgro8LD6utv99VB5+fb1QLSaodMLKl
6RuyKDX8VxRsVL75R4lG6uAS5bFEzPBSRIrYqlpKmzdtHDyFwDlN/pElKGUHH9fgpM8ze0I+CYCn
xn4npmrdj42V6qibcx71Bn8HQN6RUozgjMAspEHniQ3ZTEp2x/7uy8oGy86hBxnec6Z7JK5RtNzz
TZdA64U8DAN9BYLuKD5C5pSMTAhNWTRB6RphToYXSPG44jGemhDrUC+p1yc/+gGRGvkPywPsMkEQ
1fVwfQX5ZqQYT3b99FcXKzdrIXEx0ADCfWRhrdDc3BcJe+LY/xRUiSie5tJtnk5Ymf2aWowKz8Yo
T+xiBMcjw8lZkFV3VSmO5P+YlsxDkOmDETVwF8pNZkgWSkNWH6Era75toTkFMg+z9ra5yc8oxo/y
7OeIAqj8ewMdBHNu8ulM0MlKwogkeSehsjZXRnREcMrymjRkYrWX/syOpDiWWdMCufjmDeev2kLL
8c07DsNrhDo6qs7k6EW4EHFmyhFkwmo/M3s/JQzHWjM5g4tbKUfz5jU1VbC2u1uqUQKpSg6V4iBI
wWWAyH8gXKNK1nTALB2+9bFCpjkIrWK6pc+Hc9dXDMZbrK9KQJK+adTad/lnUwOh7wGaApTbWRW9
Fa2UNXXqBMofahQhBpyNgN5p8KdVeL9iQdMEQyenhTTCRTZUkbXnDBV196jFo0QTw5nevduRUdS8
qsjg7UIJcwm3bVF8wbblszpYyCScHH7eGIBugJ+luJT0X2eEjlW5C595Yyh7Lqoqfm121GQJ+jvn
6kgLa88U7Du8dv5InPTSjA+4gkvcnyiCR+JCTtq/jutG93CzRg2zyj4+8ON4UYCCMHJMYCyDedj4
qvkbhE3CCoQK1/k/EAE/aXh5mW1GpcQQY2a3smp+/DBaXvHr6KVe6hWfegk8mJaRmq/TFZWO4RPm
GN7lHQTP/K+VFdxItGTq4dCeKJNsSQxwfuWpeKsnHWCBJB0hNmPTAWKBjDFq9D4NqCFPoPqFlyqX
l8+j1xvAUY2dVqBvL7w5ULISmKou7ctvAwgf/fWybYpipajnZdfy4Ad8fz/bbz/CAT0uYHztizwu
2g+SIS5reg0rV3MzGfTUpJ66MhK1FMBrNJVND+VvXjMlpQad3xxuEkDXNHwNAGP5sK6a84/VKAo5
CpcEvQU4vvMqEZyiKZYdnaHl46svO140zta4Ywl4QYCVJLIczSVWemtjR0378S6dAeNSZzLY1v6f
Zgr6APzh7s0/y7HQZgIlyDXPNSQCKjGQ0T3x3mi+bAbKd5kfunsrj/1X8Bl5mWX6y4FhJVU4uMJG
DOWpzgMoCPllHtIl16LOqV1duOo3u6gWXcepNvSISKJJJsiAYAaRybHOUQG9sRzOHFrSl9s0ofAp
lS7shFb4QkwUMWidqk2c8ZuxYLVtvUILFuX/hwsOVI7dhRWsR0/e6KZmZTQYLlMm6I+/+7EOiGsx
fsSI+cs4mxNldXt381ZsoFqZv9sntB68V4VxYPVrF/IOtyqXutaNHiTb6xn2nMOltRr39d79pAhk
6qNBhePv7UROkRw6RMRQ/8R7iZQXr6Sw82eSjhytvPpcP/ht6AHoMlV6KIX01GJEQXa23ZYYu2zu
QnIUbTtoFlkGlvo1EC/zeCN/VCnIfN5mqn4IcAM1MS9MlFvdv//5iC3Rq69V2VAlgXqoivNFHR6x
7fjKX13I6S1PMtW9MXMmhdSC/SZkRK9nT6YZLYHA4I28Gfsmx7fBS9FaP8Q+kuCg1Jw23A48qFuC
+jLNOCS8IFxclTbU+9mChqw14R/tt/KK9py6pYj/xwTJaEXa0ZE0Y2FiV7ljtKPb7Nlk28oYrY5Y
WKICJB+dn9lW8lfWoNYUtuhsOAIOZRhxz1svwf0B60nGdujVyQfZuiRyEAZiSFVD/R+13yIXL2rF
+w388S7knKNpJp8j1bHmWTYoawpjdMu9sj9JobVczIdrAPF6NoKNP7I9Hvz3aKE5v9sdwS8pIlm6
fYZzDinjt1zTTJm2LFoQALCHC3QYsmr+oq2dXEO9sNauk9ZOoni5VBAwh6qaDXVnolErBCbES6qM
v6fGe9B1si7mnkr1QmeXyxOt7UKB6xXyuk1l87vtjeq6BoZ5HmtGokOzH+WJ1tiCcJ+Ut3dQCmXz
pTE2wnxeslNwXFxAsRgtTGyZYdZpyHT6EEVKkXWLDDzgj6FWFEOCMXR8qsAdyxDeebq1VV0DPmfq
6G/CjNKhiA4dV1tDyOYYyi3JEIFpU+QTr7qts7JKq80N4rXP8vh1K6cnSGDcLA3TVedsN1XAGhZ5
DQq1IfbgaxpexkaQqhVFYO17RsroUdSeqwyHOJyy6tIAYkj/07mdL/92uqUpjYEM4j79BwDosWKb
ktlUujzjCXfV0XG5sxs1GfaLKfHilUijEjz6af4uOxZ26agaJK7icAW8XaRtk/8gur77pqQRfbON
pCZHm5Ve3kdvPsCnc4fsoK3Yi+safjub5uE/eszLQGXcbtOTxBFigomjO4F4gNXxlezlKVwX2aqM
wXABn1HyGsm+GO4NdKuyRC0D9tF7T3Fza/bokg1F4k2iN+RQojFbNLlVWNJpaC53fk7a/IB5VjyZ
43O7dhDl+6aDOg++LZXzRdd78jDr84vnRYmGsffYEj6ROkLN65ETl6e6kKXJpHOEkexty1beKbLe
/TfcWk0Exuwk65Xj85+1rXeWcdUfpPrWX91XaSbFfl3WByfe8Di+WIUZwimAjyVk/jr614J0nUa6
afJm4/C/yvLPaFYmsf2+kefGZTzxmHuNV4mjHJCYyimNAPqfjeaGYkIaIHhdpNgZ6ktShbm+wSi7
WzpV1b4vVBd5pLKLrGVjwTeOc1B1094PxOtPhh1MZkuCvVSZCmnqqEpWBTfZ3GzC7RbWG6g1Xqx8
hwNIql5YTCv185uQA0KrQfP+hxZg1e6q2VX404c0IliuH/tYe33Whywt/UjDwCiP3VyNUpEDG1Si
5H3tEFE1Jzt/Y7AZv5top/nM4LceFqNtnKKo6d0Etzxk75gdwWRiF7Hi8Nco73YYy1V8KeMHYwzU
aNdRHG8Y5dQTKYv1Ie42A9zLXQVHZICRh6i4mb2qGJ+FObGsENIrtRRH1HsqPCnECSWPgtr3MVVE
AprBlXRBQZ7QfxLF5Odj0t+jqngs9FmgVXTQUvXvTzvIvmumtrqkCYIRIXW6Mnyk1HL4RrO5ZUxr
74t8z8t6h2k0BXfqE2Ce4XdNVt/cCEA+qrVscoF5f3zQXcaKbZc0QXN1wPb1NJ4b3ZWLD2y4cCEq
DE4Z/gcEW+ZjPVRSinEZ5X1p8a8cHhW7NjRx4NgzVNVZtM67w2fsgOBx287bDTsmIdGomOXDbNoS
Q7yLrSdr2a2BjTtVIPQsaOgMMQeHeBnEdpySeAke8GbDeISLyL01PrAxD0ZzORkDobHjT17jTaTe
MyJWWWd0rhUoaAhcIr5BSS5pv08pNTMMvwF1jopIbcn/oJta6x01Ubo5pWFIiSmIAeQHky2ct6Br
rso8eX2JD/UkEMW9hXpENvHCCBvYsrphzIFUF2n87rgOmEBlEGs4zYqoSyLgtg121QdIAGNFjZD+
O7TiMowVeFSvH96VXSoCapMFpwtxWOjBPj/991/wN9fMMxgoPg609tWNhVHUxKPwzwHEHf6NuQl/
JwPyh70bjor6nIBG//YGl6mNtRUWTDLRwqIdbKz0k1s3alibDhNxJTQqJncFU2IrJvlLwoWrSvOg
kPIqVG9K+80jnpo6PpAUYu0IW8BJanDIGZSqf4harQ3ScHbOBVCXmSMbFxXTGhxlu+KRSRWGdYmU
2NPNuNHLw+uuFfK23Vd+tpqQ7RT5QlvPPVBF/Cufe4rpWJe3vOLGNmSaDcYeC9904EmrV8/Tlz1W
DwQ51MOeg6gt0KsDBW/VD/oWp+vwnfRnBtXZszWHDPH3yRnDLqCpcCzoiSJvosTAzO3GrkNxq+If
UUN/oToH1yKd8TyN0jx+fPp2wajLYBFBwQ8jMW/LDqnXggLDik68ZrYLGtLAWPmjTkdlc3bxhMGw
Qfao4ixR7GcQ1zzVavZwQ3SKMPcNptIFmRQ+AzKVVklZyIMuBowPl2TI64Z0BJ2tzxh5gK9zwFjR
YwewdVFFMtIw78Uo/Puat7YGrjtbfjDbBK4SDMVJhX6rbSak/8lGA8cVmjdws+KPzVADZdyXb9sK
WdxHe28lkFlXaNqpGWhc+bxRGWiR1xq34llqV4G5mvTngMLl9qv1V5TvACOlGApHrXic3m0ibesD
C2xvwSWnIYBuJ6fUNthrqTadjQdxrXcO3b6bHVbyEeQusyEHBqhX+N0mJsCGxUzJxC7hvp1ja2G2
fsl0nLXGVre9r+twHe12BEJ1MK+vts/dkj7sdcEy5u+KxcoK4pbbUgZ1lrYTQut6IK7n80RfjLdz
gk3LgbXpqigl8AX2ucWh5aQ5Bl/1H1SDecX+J7nJ99uRk0qrJ8OkvtAetRROYET80QvPCCGKdcWG
L2YQlQnLOOt3uy4Z7fIUX4f3tc7e/L78OI6vBfAR0zx0sC2vWoAiUoahx/umLLT0IgFF7WQmwwAH
HDnCja2Hy6J8TAKrYhmeywteHrZnpekgFoDULvWv9o5J9VbNs2c7XdwD0/Gc7SwU3cwHU0Tzeknd
rOGFeJWD7Ijd4gcIvR1fdgcOTIso02y8J+7cW2ZzU4UYZwhVFfN3YtJLaZ1iNgI9I9gKjHIH1HB5
dcPte8PG9EQRPDBN6S/ycT3g220WzyLOL/oeHnzpFqTUMig1m4vtuS1HBbNdE5vl7jkWS3Qz0RyE
416N5VN3KbNmJioLMs2ZSjtyBVUHEKiUVe5A9zHcUXUyIELEEygBjGWbGg3G8Ndcc6T2j7jAlcYW
7zPvAFujd959BEFbTHieG1hgXhoficnCeFoq3hff4Zn6ngqYio41ygxVfg0oFV2qMTwgjuMnY6uN
KhtRJpqpPMqm7YetYRQcNJBL/UR8eHIdIFYWiFNrhjCukUcCK2H54IMzY5ZivRGcbBCbMfNHSfJC
WXQrUi10dIY82d1GAHIlUg3mo1uXVIrrB2RekjQZk39tw5MLGRYN2nxfneklNM3IlJBKGhCl1UEg
YBQ5l/IKMMISKCDi0XUNLGK29O00tcztm5ZYd6Ggw3NPvSDLsRFUi+htJD9FffSbHnIWtgxvSuOD
U9XiFsuND3JIdZ+9tbUvuXwOvpM/Wz84hV3PJkHYsDqJXH7FKfiZompqzaJ2iZs7QyZsnQ8M3NwV
Gl/egfvyE1/nO9SR2Ta4/qdhj32iPBMIwOegvOUSlvpjUyYeQQVHgzVWgaFGZVzhPe5UNZv5drad
HnCMq801MOqcXtgW4Sdyhm8a0D9E1jAc8vYa5ii20U3+SByPpYdy6Ae56RitAlYnb4lOiaKCpj5b
SAaMkJRu9eDhTT+VULwzfrLTqN//HQXmhlhJh2UZu9uBWcUWYhf6azuZSEaxxQBv3HecejyBBXNS
Dh8oUANJHdjDLpNlqOr3j+Zf6/xjZ163nsWrT4AUxyvDLZcQoyBCZA7yRVObaVABKaR/Y7qIC7VH
IleisFTZsj3N6XYTR/2QI29jB+j7D0pHeVoh5i9Aq2XMCzxgge4kAwHGv+EzKoHObgcw8Ol6Aeb/
yaViqiCy+fOZwFWln7Lg+DQ0sk8eabi1UOEOfSbEokPAcFhCm09dTEThwJ4JKdCkhxWkGbhzTNIn
lvdwkquWLuWrx7uA4lyhmaBNXz5kRTWYNJ6m8/tblDfIdozAZEqBTaubW8Qe8D8Qqqt3AP8ZQDr1
SSiKUfPge4SWKkNU7DvbosJHuM6Q5IKbBU/YYOetQ2SzzhQf2VbcdNIJgVDh2wBZ/AbRqnhfWTHz
eSBd0v3GrKs+DmLMrBQDwZeSBiqq6xwED0gMtIz8PWK0Iwo6spC8O42ECJhTX88OH2PEENsj1hkZ
+SCEIrJA3xjPZSFdKrASHctjdD0mcthxc6QS3MDrj7I6LIv6yhjTduV2X50qbDVY0qfAgx4EeRL1
O+xAKBXpYCZphf2JUmXBVVQmsBb8bGb5Tiq0DqEm2quv7a9ooNUlFCnnLFnvyMmZ9hpmDAOSFoQ7
3Uu7LgVgmDoj44kkdV8qTm9Je077uAD+DPdVCrQUscycucR/3ZdZTmlFuL0zCED8FVM4wnjgbi/P
qpMS1FQcwV9cX8z62ucyiM6JUC89BuTjLzEX/xJ07xBqVtQebXG5sIfbNmqopiTimsEZN3hoE0lJ
BmUC4vAbHETgqCo6Tjc6aPq4JLUatCqvo1yeYJ1HqQklT/do3Q564Jpzet3uEwHo0rtoAa5T5z+x
voitpiyWsI7BdbLaZuqyRVQ5MkBbhyxtLFRapS7IqlNuuGehqfJ/R5Cz0H+RlrHNk8Q5uDd0Sxfd
/L4ESAxWDWYn7tQ7ZI6PSQMjm9E9vLoh3SvfJqISxjoka3kINScFaimuyRIAgiN1lYNtzzf3vfdX
Hor5C+J3YwXNJRdF1TGqRJQ8ZkwDuDoSyRY9OHKoXAmpuyM1uZ0oMtBfV9FnwqDwRy/7qUNh6m23
WVynUTR5oRIwkXOjSP1fC01yuY7vCAfOkgipYv25F4T0UTmkXeQyiTjFog6eI1CVrDMeXEjWGQ6g
0yzfOiIdNP++cFgihPGM1QYpjwj4sPQLPhOkSibaQqKX7WAToFw9+npc6dc3beURTKscpXRQVBmt
QnuK8GUVoPGfVb++74rvvfNbLYcwmT7or5GU965ui1jY4gOnb3UKz0fqqyLWzxRHqEqabtW4K9on
mYIXKB4W3wNFT62CG0rtWqelM4DFoWGRSi1GHcAWpgY/iAjrGShp2F9TxisJFXIEZ2ivdRWbPlgW
cLF+s2+cqnkZRNpGeLL+dvWag2dhQcyTt1AgTZ8X+8gMBUyLXly7Ya7KlX4NJTGIZnYrHI1Mz4e8
dgJFlWyLu3iUnGUxvc0WmDhMkWNn6t1t6tSkEOTzMF9r8I0bFVB49ZApCNCfmzhKCqTJUR/pFEQd
OJFaiEg3CNt1R0BokF9RFs+E0fOgyWimwvCoUGfpuunr/XbkXtpKPBfQQB+CqjrFRjSMfOU8hfNG
nsrscbDXt10Kr6DymLC0ujmyh4BMr2INh9Uvr+K0dmjlju6x/otoZyhLuqfnUbesxI0CjTQ2tlEq
knnLunYfUahZUdqwlg3Pw7F4pUQG8VVNpe8blVNOrgf5hSZuqm6oDkzV7mQQjusLZWp+xqJu+Jtd
8jNsEBbEwY/kO493yB+7p7beDBmJQNztx0Bnk2M5hPNAPn0av3878YjgwEiQNG6nc8UV10vxv2G6
GJoz4eJdRMtGHSe6Qo/StuySHXsIeu+6wof8G4gCgegGZ8rx5vRulA0rQGSxbWlmawPeWnUCUu3A
2FUkGZ++JEMM0Va2RnS0AG1DMo3YeS62WMrpe4qLJbEjJ4/xa4zBBRJokYk/krbkg8ih3bBzUm0t
RkNmrsE2kV753YVJZU7+4z/KEAGDOQPQkjXtCKZhscxKTY58DI3572sffKhLd6vABs+SSFY8f5cw
9KxJI0och7F/6lZPfgFJf8UaHqPa+SnWlTkJo3NVK0d+AZLN5WWnYvTBQZL/arpfehsu7pqE14Rl
gfTB+vO+oqfPM1h8KKZc6duAeA6IFyf8IB7kzte+jz5VXoKYBsrqLOYFiGvsEaDoDY3FmXNG+Y8b
tY0eptgWs3Ulhuq6i32V2Xrd7rGi1nnZ5JEd3obVcGTKtj2fNuspkx+q9XG4oQm6o/gj8DgkKmpN
gVK6jLd42nitKYBObj4/KTVnkMh2Tk5ZRs4ZAltCdOUVlIUustEEep/t4oyRir5MVubugbZOZL3i
Tx4Q0iYQ/PsSG+LHOSBDDtQPEYX+a1bQAuyPye8FdJ0oG9VosxHYF2PIZr50N/UYTgeK37Sm0LHq
6N/KP2BPaGzLys0eS86rgp1wkbbnPy+gWm6JBn1229jX2rapzJWHvbVm6ATVJJTBM3083Kb2BVtN
u99OXI2UZumHOe7EN+K5kcwPjS7UUNR3mp7jgH3BXLdJU8iXHWM2tq2SRvvrHCaLpw9K3EXDvB9E
//hOud569eWPCWomU2YAWVArvGDO7adkTwCYeLIYK5cofkQ1FyqfHwQ1kjNQ40jUsFnYMu8Ffj0U
vpUVvkAXqw9E03efkw+Qcnp1KCmQ0ksp/ZmenFFAv7M29m806pyIjJJUWvGxOjyvMOuoGw/ocCfi
qTMuD4IqnT+bRM5Xo1hotqdwJ2RtKIJqKtmjlyvriLNmHNP1g4I5yWf/qdPNsneizh+QAc86AzaS
UOKt4gYwKPd6hhF9j1/3UPavXeFuefQ1OIEVMMrGEEjVk2WSGwcngks0oZHmJkMfgTR1yP9sLce+
GmkdUEPHbaN6XUpPzhV6w5YRjvqAATo+0uelX9wQStJEj+wt7IPF6XSvLhLM4x/FLjtKqEETX8LQ
Y70uUroRKMZVtVExiX4nwxGIvV9UnS2lrCZ4Xfu5FfoKzeeCEX4QeFwjLtug1ztxAg5iiGF264j4
ZrRUmq/Jp1ByTagrbWZNRxhr839tYDPQU6GRd3VerPPern7ix7sZ9rdbxqJIpdXVs7jFPncx0gjl
MuUsYBCPbqi4SEBFl49Q0u2xD94BjGb53XqlNYN2jrc7bR32OiRC6bAIF+O6cEAt7A8/6u5/UZAF
fNEF7eF8PKh6Qvg0dbG4iYPh/dcgadeF55OPB2fBQzv/mu3oP3d9nUX4QyPWpkMJxnak1BNeZv+u
vMYsK7Wp+VEd5xOpHjbZl7OdT9yOZB6H4pVPQ6GD5CDgL/r2pKlYN8w5DDW5bGrDdudoiJc+bHsE
/hou96xZj+MrJ/meDR1/7Ml7jUkBpSXZ48KzYcZxhQZHeYpSbmoMkFNaryuOchdQmU/zVRTzvCex
yLtAtmO6U+rLQyDgRvv+XavKzJ4QoKnXCFL59dmQRVU8REfHxe8V8BSBsSrQ3qSCo3ud0d5oLobz
Ii1UIepa+SQxYOyAKxN55gg9elWa5h6EeY/irMAQDa27ux+xK8UMawTqFz0x2itN4R3UzE9eYvFw
ch7q3Qz5xo5mNgPbH3qEFJ/ciK5hYlXZmzLyaCJQTgaSilMo7LdFmafFy45FmCgM07RW4uPBxeru
X71l3X8vqWn9J1/uo0RdPOf3fgMADtDPZXvkCg1Z8H2Q0AsJgcJTFoSi085ZV9A7G07GGcG7/LyX
P4s5osaWTrHr1rB7iNpmfmIP907meYyx826IUj1qpxb/u8YyEOZIy5LWKQlCWKePpNIrg0oeJZ6X
WMotlh4XNXaBe/hqNWqxbksLp7HL1P9dZs50QLZFos4ws0KI+Rn/v9swZkUT3zRqmx4tQAcpQXn2
WGIAxOtIB5Z+1iFqY7H2WXIPfD8zCeJu0LCzHcBaI8LiUDHnECusVq6CkWyPx2kh0tcyG1ENyPnt
gCT+sSHoVLWs7NuLsuxw8/m9TtOZdoDHVufI0TpYmMC45KHVSUmNw3hNJlPQqD14ex7k+hlZ09PO
fl27XrfDTAyZaXbmGYJAgP7hWcbMZaDrXVegK8Op9MakzuS3Ha/eYCOnCVXDe6gM/mBy38aT3CuS
+aS+g8X6/sQw17kYFPwQ175ALbLX2WEurB3qJkBUTcvCis4cdBm3lmPkthJ1bkU4R23AO99v3XXo
wX8iu74sOkeGBXfKLsyHNUm7qp+MTlwIAm03cE6WsGwdk8B06KHVnzD+oPpnm6orWiW0c2fFFeQD
AZELZF9Yy48CPB5muMld33Ek7kMPKG8ukppvqU0QPcZ6ZGDo8cP7FvKvwMd9+GJQuFYHZYEU7DI+
PquU0u4cPvbAzEE4aDQeWB5bKnOdHR9Ei9iyRNsRYMuLeHrQ/NZimACzHa2VxPiWo9F0zK/4WhrW
vzNWfEy5yJKfkKkUISR/oBgknY9OA9XIaa38wuG5mwfR5WAVQCE6PStG+eUw5GvSeokVY1i/dBdH
xU6skb5oOUAp7K5xhVeZ5qJuLOklgT0Hvl5Iz8IMFfkg2sIYTaM9N7pjWZ1W5u88TM3eTENfapOp
KahBNNlBVCFqCnnQnC3+ki4NvZJeJgv0A5/z0uDUyFkeqXo1B3h/DVS8VDzr4U0l8yxr3kKYp05N
mwVdVptvPIEKxT+dS+nlSeZXg18wst6hiRNN9VtV+dTKoSgSuw/4yjhyUV7D8ljuJKAde8Zrqr6R
C/Job5wfQ3aiHSkWopq6HG6f4N3kKNl1bVrN7i3d0KYNQxa3IwdNYGMRovmepTFUTwJsdA8uB6Bi
SVgj81f/9vrMvBrRhWmEq9J/rxQAdrFx4fV8O4EjySanYbNgNaQcWPBORSSjJ/RveXskTlsD4JJt
vEz+wfAzRyl7+6UbP2/hJA9KfqaQCizubkg0BDGjBBiRzCopShwe1MhYafKa/WtcEOp4LmTPorez
AFSLzwxYY+Pu68FJm0sYhdGisBQykokKNtjV3pWYtbPz/2kWmfA6nVjs/dglFmjSo3mlReqGVSio
xDrB1NSwWQ8w2oD+p4rbPlVstdC6rPBLKlaAFewLec4I5R8eUSHG+/ojx32LLRaV8wg3GQzTEzjF
P5xOKi1zzFRUTHYuBLxEUJmKYsY//fTMc4k2ioV6Bw3UG47/GDOjKll1R8mTkKFBgsEFzvL85jgR
V9DPjvg5Cgtqrr8XbN985nXcTRvuZxj0ayWgTppdz2tobGxO2Q6Aon5d6AoFstcr/aNSo1y1mwah
AKAZ5AZdCZEJZSCSXXF8cU95VjeM2qkK3Kk8owCeL3L3+TTlpfM30wxB3pBKOicENCY4VPdnYWI+
I4cgroN2YXU/DJh4wFlW5bS0agceUPzeJC3ATtSVDQG1dQXJrOcbJy4Fd+tq9tGh2hM/bU1GWnr3
Uf5SE83C+kLqm+xPrthffR3b2xJkiHJQoihUTNpULAygAGpDLVb4mefP8B1AXT0rKh7aBMCItHij
ECfp3a7Y96bMECddhCof8jxbxMxR1gxtvY4/AkPfv3/gHurghAB3dJvcdNBnQEwrhnglX/n6p7YU
2gZ7oZJc8LMn7PI4fbYSF1FSAWp+zQPqdVdgn4PtrMd0zNvmpiWks3CWvsm9fm1Zg675DHTgEbGr
8nTBXOfUFyN1Qt6fW294ZQrzAIUEHMokBGQEoAnyG/0ZCpm9cxpoUEGnZ7Y18ygcwmk7QWg5X2NA
D7d4f+PfREllo89XIz+mTyRlyKKOewnHFjz1DE7m9+n7JpB0Kneuq5VSzg8Yf6YXjUts9eM1981K
pDYKuTjrv+z8baWw3c1tdOhCkVbGY+Vgf1XmbB8zM0K9cujfi+ppEaGlrcA+41289Ww7uzXe7QMq
SMiWkcx55RUIDJznADuCq03RwVHkCHrxsYO1Sfrymmc2kT2fcCZ2i/fa55bSrhDn4SLoDsgXMjEm
8leT3eX08g+njv+s6b+RJmSBTiCLaDnxPUxYqTqWu8EUA1Y9bk40j+KAwJQP5kc7tgnz6AFS6QUR
ewks6T9ZBdcbi6A3hVzP78scLyhTEIhZMPi/fEzE0AKdqkaBoA3xX1ecpFUPOLeNNURUbc7UjVF6
7zLXWGzCqCzJAuLa0ineXM6pC6gCq0dvIsZScle4euVRXwZ7ePOvUbu1gsKIVMXkoVuRmrpMIuXo
sTw4KKjscPw84iNOhe98c5Jt7EX83HGAHHe6CawQr4SwemIwV01/JQ0mAozD4ZUBN1cVig9iL3uu
/yBQowje1g6Xa92LM9pYIzpdRclZosL2nEKcG/qFnpEf6S5ba9FJ7gyVFgHD3oXN2ErSoun7nPuy
qCxTrVA83uW9ly6ykTRKaA0VbkfWk1G6Zp8YMtXFXkTolRXUuersh9RDz02Rv2wOdVPF3Gy6E6X4
wfZ3do+4GfcaGbzg2rkOj70Vt8lmTJpWZm9tMZ+7QxJtrgD93/00XTHIWk4vf7/RJLNsPWClKyX3
rGKzBCiQtiq805pHSpF3vjwCPEyL32rl6nTkb9Tvmqu+6ZcRDAPMLObYVQVQvkXxvAHo7HsC06W/
wPVZZ48TSAmkP/qaeb+a2tB73Y6/oX8GcB+CrYyiXZ0yeZ+cH2q7eu/2WJ6yq1fxOD4CvrUSqrZc
1pHjUJ3U3cEkFQKfkWWI7eNB7LtZml1X2tTkYgR6/D+Yr41be+vN3uVArzFgugi7V7ydJX4vxGnV
DGHX2NTOfwS1f9BSwahdKqDB806oJYoKq78/pnrFhBYVJeUHeef7rBbcCfoIry1a7Gm9yoCaajrw
YZiEVT148wjRFk7wFyH13Syyxi5qvGwBjpt6TJzCAbEGh9Je0SUHLjszZVPoL7DmeUvaV4TdWRL/
a2y3gBRHCmb9hfPHnCB/S3N15z2BbYHmVI3JcIEPeULeAjpsFVjDn+NOhwwzbB7fv/NKF5jT/GZq
gbTa9gsOiKnGsiNP3UPjBcAxTmXlM2lT4vtUGKSoFdebXWAB+xOype5KfC4+T+3c67w6a10Yto6L
cZw+nOrhhmY+0SINw84lMTVUTQPDqop6Lxzfh4PIMQeECMhWe3pjaWHDB7ehyMbEAxCyOyDiOc/w
GI7t/Eaqw4srjkrBEV8mEudDkeuX/8uWfyvNefEVYrMy5Cbs8nj/2wEA+iFf/371KrHM2pAsGp/w
X7JV3KbRuq0vpiqXE49GOjqQFAvMmrq/J6xqrPSFvOzphb2UPqsF90Lx+T9gXxhG0LqQcSadd/8E
wc+Z0m3IBVQFP4LbEaLdMCXmcdopLv5lZUyGjLzBb6N43cXVE0p88MEL+Hk8HpqlnYlHwIJgK0VJ
AfoPIAYi3O11Uoh7iHiRnkJ3CQ4fhX9hwtZxVmzTfQx955sfD6E4jStlSTdaeU/MLZAjjOEx/J0Q
ft2zTgdXwlAMwjclLKk3K2R4WyAkQgY//Ujge+wMaeK1NxEQr+vy4oNs2HUOgm0XAyc/8JWvw5oA
41hys+rfer7XvIbspdP5pTYlPT3BX12MGz9/OfEambkhL3xuIKXWKeY9STLUv1Px2PqmrnsAbAKc
JplrAG9exU1OWR/Rif2eMQciYhBG/z+2EtAufILdM4t/wz43MQbHbWpF3z+txJLik7UVaVMF3G1l
/6apMGLulmeyhknqx2SA98dLXYF8MRU6ZK88D2ojo6TIhbE/gd9F1bgYLS4dANk/z/fwDBw3cl/K
8BxAPEbxPK7RRmu5T+3lOCCMimJlPr+7grnYfZUVOvTScH9va5oJJ3tTO8a8qRSi6WTNNgk4BOu5
kQ7aqaiOXV1NBRyr7bgXgsF/7oKmFrA8iNCf+S9SzCjtoQtDyzQxZax+ZTU+l1UuD/e2GoC4qhpV
b9/Rj8R2xj1eEM/ZgN+qONPhWcnPWvypNznBqQFM0ilGKg37oM0B0IL4oNdbxeVaZ3X7/1DIHcj7
SIWRX6KXALuDInWSJuQfqISx63jc0rLcVlT8vYxwAbh2PyCdydrSYss8h1dgWhtZhYTqqVd0+tUK
PjavsBPOY2u28l0IXx18wN6yvmXLycPHdAPpN4Dzb5zOoHrP7g0Fx8JbwGBhrOUySg8RM/kH2iTa
HpeLDAwyxvSCx0ucZTRbDfdWCCAv1XJlx3EDWLP07RwXX8uZe5bUIus1HZpy0IhHip45dl1HlL57
OpCjb4+8AzZ9lf0A/Nj2wD7i49CchxTiEqcOdkJ934pNKz1fI3MLI+jo7bfw7VCvhP1G6E1sUy9U
+CXYzwDVdszI2n1H5cb79zEajPzaf69oNu2UiPOIHH6HukNKbDoKgRoNS3bGI44T0IBEdeQErK8B
/KIJID/nVITxnkPQirRU7gMwA9JixLxzP4goDePVm9jv6PH5dM/Cv0X0morL3amNcKIbi4icfJXS
7+gkmYISJq4sTFL1JffWsCsPii+XcSVHJQy3ltFwmMv/D6O/5J/4/6WHABaSpd0B6/X78n047c71
xw3xucBWvTqudqVEcDSeYOuFJAv+716VLlHwKWhkYZWRvKh5hgYlxgj/FrdCuWxQTdrcr8MFy724
f4FUJ4JfAb7d0/Bekxv89yi8ZlVkdHFY1VQpEkSZAnYk1SAILT5JePk3n2xVogFCrIBONy7ThvcF
TE79ak/K05bw4vxb2jQoRmFkWJAo665yreKTwNK/J2hIH8C3Eyq/ojqx0DbzN90O8P00RGVhYAPs
wLxdzd9u2NIbXsuQQiZba7JVf6JwAVSoUSOSYrCdvoCW3gi2MaZ+0EJAwRhvj9DHrdGcNTDv3FNX
4yUQN4wFtWdtEY8BOdo6kpAoAXQpgoDl/u6lQhtKMZeLZ438mbTXbZAdaFdFDkx12G1TqZ2elgaW
aRcD/lnBxgfKbTgxhQITSK3Yjwg5c0HEU+cjE7o+JKfd3TAUrAiDwEjfOde4UzCaU6GnedCKdkX5
U1NoDi3BFW2QSGQVe4cTUzlq7JbAfljMvW4vSnkHQrFL9ipbCuhu+cOvSlHf712X80BnLTOPjnBJ
LkTEiaxhUG4Ujyhp0oYr8R1Yr6GQX1S7TiwMLFwGvlECnBDhlk9DNDG2fsh4rnfeP2Sk1riCyL1t
3AVoPmUiA1yV6vZztcIQqgYalyjBucrmg95m9CPRXH/WVD++aPZX7yMsPk3vXjAHDTczHbfqctnD
KX72rHL9AAu55ZwAuE+01YFTRHTf0btRUyfTAjkp418zjE2pAkkvF4kTZOgZ2aoQDU0VH+fTKYHb
EdvNx1o2wtqi+WvCDA1qtrfePvAN3L8bp23AzcyLYtGyneHhIx2pBqIyKjqtepSCU962vhruOuF5
Jb35h6qMXdOyOr2jBxyHaurnlqibYyDiG8H8lB+K8OMHUH1RD8Rn7sgxCtZVcR7RnkHrHAosQCJY
xMiHCEtW1pWncgDhn+nEQzcsx72wtq/TTFzo83UH1S6/25icectY1e9kBtoozPaDzBxV4uhjKvan
hJ8uoybQqxlWf9aBhJG4tauH6vSOFmRlMn+yqKpl7JtYiU8GUAIZOW125OsKPIJS4mkv0mQk7ozK
sRv87ohKWEnrgafjHHkb7RJLcuYtSdAioFojmXy0J/FM/5Hu3+VOPnFRwn5gwyTBTUNlpdMRf6KX
x0PTdEjcKq7GfNc73b/wuVYlytDCSS/VsxfhPeoU0QhS+2bhLaUlHFUOp0VUDC+KI4mFcJP9KZwm
czKyECupx14roX//qcCEslbnUflrllyG0fMkbYi2GVFecn75KykILYAZPs+8NlZgomPrk72thMVo
FdK+3TbewcuQfugnzVpRmzIYWKxwTEyMQmcNbcEm1TboSM5a6OCxMai2HodAojgvsXRKMLxNMMcb
MyMZRIIV71vYVAoWZW4GFhnE8XlFayK5L4znofD4+OvsNz7Q1kO+wNoKNBAXt6ukTZ4anu8mgYFl
m9OIZxQyhcSkzz7mvcsYmkrFzXXXilAuSU5e3lO+SvCW6fnnBoyP6hrLd08vPqFcc02Hugm0l0Gi
U0UvEH55aWjpagYcvgsG5imSpjb+TDCMxmevO4YUH+zgkhXIJFqO/H+JBHFVqrS6hDo/Iqz5dO8L
j9B8pQJN+ilLSweiyjKRU42eiQhZdpNQn9YsMzVzxr/JWidE8b/ycYXfFuA7Fie03W1K/UzczmJ5
Nshlsce8IzWOOJXqgNCCGz+bJ8dDeJ5JAI6feGCSS4MjNiRkHLR8udh0gigTPEfRLMpKDALNc2Hm
ElhYlF3hwBzcho9CcjGsDOkHeltDVRCKsZCPIdCHuNTMkSy/yj5OKGeqiGpo6/Wzb4EftmhTAv2e
OR6MGYs85uYsnLtGJHFuNAyMY4vRZXfvrCo75Iivy4cUlJShqtBR8B1oC86xsD/X9IfZGV8aKY/O
no5hv0QrPHvK2MEGkEoxXzdn0rMDiGmT+Cog1bl5MRa47pkiLtDGJ5YlVpBkH10ZGWCxiCTZwVwA
jqm0dz230gaFJau1My2p2zER9AiE/aejRQr1xEI2TldHt8uE7SZ+FnKI3oS9xd/ojz9JgN3IND8P
xJhja60ZIGBstRujw3beXMdAVXOO5cyY0ZouOzsJfC+QYwZlPD/hBPKWZxcymESfy1xrdHiZNPKU
HOPslEatxD6abW3H3IKd8CIjQlx62Iir13Rqp3TfiS1nZDHWO86jjbyI5H2Hdf6HfV3S1DfwSdDQ
sAr2RWTPfI1q5z5eFxOKa6Qr8V+73/jti9aJG/lM4bTretoOQa+3wCAVxTEJXhUWTYXutRuTz3KF
8imZtbBpfO5SY4J0OAm55MUEYhwlyWJI2b0UC7uJty4BEONhWrT1qOVQRcxBxsUqQCnEQb1QXrGu
48+Jvqy45WQKG891ahTDxyoXc/OKYAWlHFMfob86ut93dVFFRzfvZbSVzWE1PcJJgW3+8FEt7jbm
plhL1YM/vCUtV0JQrPmk2o6Sq9KK5hWlnK3VQny33cmwsryluapzgw7jSaV6UcJkvq/flTgj8VNW
8fl5ZaV3dR3Ec9guJCN27xm6w7KFOchZB3nb6aVYE7pY1fnxpdEe4RLhJwhh140+z06Lv8cXOV/K
q5UH0TBv/dMTIosGeNt3JGVX0OVxPPSGds0nkMb7biTW/zbb173ATKfwja2td4NuPvIwcmv20rKK
T/mLIvrMcpeprV7TmagjWLdLbk/GC/xa+G+VirOsIVGXbqfKdgNc17UxFMwY4NNPko6pIv3td158
C/aFWs5XTAXL86IQ5709zN9kQxn4Hisr5zSjj3DNcQDvs6gmNaz2Rm6yGjBbzLpohKOTsw/guoqF
9MdXli7QTS9YrfcPBsqpabiNSZx+1V49Q6eKm5XIHtwYiIDSF7F+F3L5/LOOoiu/l9lN8LYNy1Q+
mqdCxdxC9FME03tVHu9Q9ro+PqJyiy6nJUuWjUIJPYegimLonXv/gYlN2jHBhjCun6glan5CpvxN
gyFqsN+6gDqLLSyt+y8/ZLV8oFmQSCZNp9g7E1meiq7lnDmb1c2I6W9T/A9UStW1fNCjz6CKaEO0
sT9CPbldBNurHOL6ontPmEW7Xc8vbz48VEvMQ46Mus+zJy6RWjfRygzmbMocjl8nBwyhoSWf326G
Bcc0d4+3bo3VZnBoNWnO+dzZ2gdGdKoeuJSIfK1tSHUyf7K1UsX57wwIvyUmJHJiu6cEOT3bcqnO
/ljqg6R9lXjTcCFYi2Muflm1atEYt04vnS3CcOrHsZCg7MWvruS6amWvJkNKyTIqqlf6fCMhzEV+
T7wiTK87BBQds2LCI2+2cf7CcOqahnKPA7a14+rCT5CDzVTq3/KC4Uuxc4DfL/7302JFhSx1O+ae
mJIs1wUHDSovSIWa6tRavy6qH1Tq4ZkGWK1BnSzpHVTzPd+hjvrsriLHEnZE6rauDzdg0/OwGRre
L8KBfKWIuzFqkwtJBdkdLOV4cATdqepfuuEzTux9ZOOgGDi0HqlwKNGMIATyAXuwDDeDAGhGl33e
8Mh6PwiyJ8o2PxLWUWMcX+DN7k4cZy1kISA+RnINW+2w/0WQ4Jeu+rM4O6o8OS5L27yMjr9cw3iY
bVzEELGjnz1sKXmYRz0qx5zxf1FPl8onN2pWA+VImKJTghlnVyIPKybim2rM+kvcZsfrqyZnVJMC
sD3W66l8MP52A6Tej0U2WkWhhcWvt4v+wG9Oy2+EjmGHriFPmirb+uxPblPTkTh/yXZjg4cwHwNu
X0ujLftwsnfr7KmtMqEG/R50T9x3DsxfSXWQtTcjg+frU4TR0HSHSDXMvvdg8yg+ayj+mZ/t24x/
Omfbuf77jC1pI6e41o+b6mr9/Xvxu3o5Rf6TwkW0EyJrhkt+bWtBKGw0GuvXiLzIZsF7hgO8WJ9T
kYfuuZP865bSZtHSPnV7BR/MZsIhKq3+q/Xu11KsmNyK0lbw8VX/V+mIM7V3PvJd9UR8Ich297nn
ZNpjQppCuBsZ+yXDMlxfY5tkMngG3htC4t3yHDET9zyPUJVByq6z9W+MWFoAWRlToirZ9NIf3DUV
LW/zMwmkW+u+/Ej4Zv0T2jxLbjl/j0zKJP8XhlliIg3w7F9rtx5g0O3ALQVDwDH35nmX/bByo318
s9fi3TlfBvkzZXDhd+m02JZTtZ/JDlYUZk65FhdECmxlsCVVo5Q+HCYRlOXDHU6y/h6SRzYUBlwT
btvyv4YHYuLS0GGTTDts9fJigRkw8BphwOz0NjXDedYCgvV8pURogpSC40Znb0ZRpLMPlFWFXySG
KWQmAJLO95o5D48SPBAXtKa9TKzoZqSy9pGzhXLMmnVAo4QnjAfsIGSIimhjBkcP1UHju8DzMWgA
yNERUHtUBmCjxt0AYXwMRFIiQUtAX3U0pZLZ7n+k1hWQHl3fFs/juFaUG+fMQFkvKkg7VDEcRdov
dOUbyODtbNNphmXD+9eDQOnwaHmks/D+R/wzQPdXCOPLqgErGw+8hjj4hMuG2PY5tCI9uERVGTCs
2PQd9F8Ey4+OpRJEgpRvsL2Ylq8P1Woj5QmvBHQa7GTU9IAizpBqu0dm5MZB4moo08i4p/wFrcbV
suy6WidifTfXK/UFPMlE0w+eMKh6zfBBkex6qqfLamJVayvpWlbRp+JWgQQ5DOIJk2pFGnxIOCGx
0p1q4TE369pj4xf8ZoB8XVv/Ec2RIWebB/nOZTkmz4sSTTzwTi5tlfzCj/Lw0/nELix5qRr6m1va
m0CFo9Jwk8Q49OVUWrLIrXAyBSgA1oqedgPpCLXOVtR/EiPCix2XyM7Fg/o+ypHFIqR8emXtrOBa
+n4AVfEjrUKV9GVKDWnGLncf2NoE1nUgd3q89O+tWudTZSqT9bAzn8Btu8KwBb9oI0o5DMaSfRlY
CucDYXIrz2JM0lQ1/vCdTQ7s6ER62XPlVF8r7Nn+6iVuruRcfO+wvanxcZYh79pLLNqAc5PZ983g
oRc9jiZ5GRYUlz0a5oimQ1LzyEojkYAt18L9X0EeKKYIIefGJtpR0FeSd/RdufGKBEWxPz82G8BZ
yn4CdrVLxqtqMwCpR8OsAk59YXTk8KO7Lr1oFdxOO2mKvDOxQdKI9hvy2jS/D69sraRenejyPHQ4
0QiB34FEj2QhkaD5A5cBudqM5oB12SRxpr+IPD/qBlwojyVHRnZUjHWdOl2c7JyxjqxNjFIC/JPw
7CvWyDRHixNo1F4y6XkwGoKrrDrRBG3Uc/FbZDadQkY9mXQkOg1CYmgVKxCDmzJYxkltdhsDgLji
swyCHKZ91J/ic2GscFV+DkTPgjJpinYxkuf8D0Wa1iuHmSBXF/L+yHm05dB903Me7nmxCYLv+c0H
J1K94va4m7KHpKN3F3U1jstLqMg6idNOcWJoKXM6nH4gDAqwmz9dFFXqm7oc+yUxJy66zgcF7Gtk
GHoqyloxB1/1n86yAUnQmnqmNw12RHeQp6xFwMCIvgKGGM2pfA7IfcSLwhEy4D0+6TcFr8O3ScqJ
4SZTRSfG5odG9cVfKBsNqO55Yh9+7rrzDGfb/cFaobhEO05UPLdg8DjFLmd/9KW8iKya+NLv4uJi
joN7xTzWOBrt0Q9vl5tkz0bM/zAf9fb21Sx4EENu3k1pkj7ZnIffj9IGVrTTbk+g+b3ULv5WVbJw
lDYMdmcvpp26Dbt5LGs+xmlfAeyJBG2Ihb7+6AFP1mb55288sqE5iub5+W4qY4qUoro7hkfUElRD
4JhBoWdYeXcK2Mct+TAuAQo1lDQzJ9eItnPwj9DJVOSXfVMFKqCh37kidzRT/0BkltZq/qWd8dh3
HJvb2M/6MUWGSWTTqBKXdJVUeWeNNM5hooBHUcdGrm3QaW3E95AS0WjCK1T/2gQy/+sMF1VK6gtB
lVlYgZvPBAllYrelmRSrm+ciy9gArYEbPsRRPXTzEYsIX3U4fDFx7xoUGQiEpzNyTShbDUtcWBAj
eLa2kLDs/p3SI2H5Ra2tyK+tzmd5oCWogRi5K+GCHiPOBIXNDcZCN/Izow9KCpqewW9YezxaxC8z
W4nc7TBNEksccKdZZ0Iv5V/kYTCXcqxYZP01YkNA42+01wa97q/rDwwDdU3HkS+D+kTUgN4VNdZu
8mCMGpkS3yVWdVTlLDWW33teNIPCNmkuzZPPgHb8lVPR5TY9clYlbhvaP16UcreuGuVqdPBnJ0sz
pUPyEC0/cK90BBQe81gUqQK0prBYHXlBTgOIzoJ3767tTqtps+YbK9mSm9A6qmMS6edzzS/3ld9E
UVDNMJvJV7klQSVK/bjJEqev7TCKb0VUlhoTqL5KcziOCrOJUKGyDi4BBgjiHTTmb6Sf4FyrloBC
qZqHzL6D3BYQH4cnq4c8KM9YyVnXr+EAUSujvxht6A/Fzd5Dzcl8M7Y0fcSImhCHsp8zwUrOQR3F
howcfwE0SG9JVoEW4bFC8ptwz6Qp7+Udx9SKMqywktwRo5d4Ps3zSohTUJEzWDfmyoaA26GZ4De1
yfUjOxiAa0fE8pe+lbkvJwRc+H3kaldRzelpIqQ0U20xUNkdhYQyauHwCFQvEUsZBJxdLFPY8Zzp
WP9bBBiFwLyO4ybL5+5O5pWfAu6kVDOSCkSfjz8xf859n+D1EiIfB5qcGTkAvXgMU/UNCEsDH4Xv
TyIQDMJwGAmhgqrSUmmQgkxGrBvMZ9X68ts+sFJohfWrwpzUWg52ODxQGMnOEnQmyhRiO5E0GHuS
QCkGQKHSphIaeG7q072EGjbSMFBzRBeObFnP7VCWGvB/xGmVXXlHPTl5CmP+NH+/Ule8K5yxkRK0
M62gywQLvEW9b/vs77dL4j/I5JRnWG3HzyAt0Bftzs1g7nhr0U1btvY+/64giJ4IE9d+829Ichny
a2sKiaq7GdCABAcgu3dCgnTET2nIgi8Bi8u1c0w5T4eHvfe+NV70PskWP32MnaxbW64quhXiVwK1
TA1kNwKpWE8gy7lWn4EHWRdSpDKuhrYyn9Tde/UpRNSoOhHCbxP/z/uDUqC2YnvFCv8FZYkh5FLQ
4qbFMFpKWB6ehkM8nzPYdw7xZclF3ZgJc9r3Dg8NKkjTOJOAQqrrAQglFUu1YkuqqpaeornCDdD5
2BOfjO7BlJ3mDvXBdHEwi2vMwLDLx7btrW3ry7RHMru7ZfV8xtZsn682cW1v64FP7NW3iNPEDP1P
Omo9XN6pVQree0HiSKPKuiiO7fkKj6ZIy8i+cZq8HtZJumBDqV7bghZVd0ev16AwNJu79Scg7oQE
OGky8u+khHfOdiJC52HL0Y2ob23dOgBRdbnBM4XSjZZr3/3ECvJ+1Hjt1JGe4HN45ghRlqHcfiuY
jLjQo3ajjNXhKxXqND2MbN/St/VeNS5w9QpRWJj5aVM92fZO6oJK1Ck3uqvk3GjMm51g28uVFM7Y
FSSSb+tZLssgKusHJsrmt++LpdcTSvOIXRReR0yTq0JMnpwDgDeEYf96G0OITUhYg805RxyIjKv0
q86LgIoAsRAKu0OsWvC8WvxzVDtnrxyhOB0ERI+ZYVuO2RbAZXWXAaGhpe2lqZJdpqB3bbuIMx+X
lbK7CwbeU5FSxuTi4gNDq2W62Yrt6gKS4c4FeRibMJDsOSAP9HhGYO/nxdI3eJcD+GfyFTIbaICY
QJ7Qd4DiGIUW+5OCnpU0v6ELDmsX/qaL8937Bw01j8tGbvoNTT7oYGxcubrVXHPKt1TsiOYDFcEC
rCKDnZPh9Wi8whaN6lXKzniEz3bhIYcofqL4aDKUJVy2918PWIaNCbeYS4RSvu24QxfIBo9KadjJ
1Ix62O/gqp0Im9rgMvcyDyhCvJ/zZt5zz8pilRVY6ezF/Ait/PKyieHUflrfpVEs2t2/3nbr9mwc
+QPEvmgFz5eBCIy334sh+bvwpAC2uT1/1u/F+5SyGJEkmF7yy0YUNBIETBoIpBB1VJAbl5qVuupL
VVUmnagYZ9NP0E7vOxW8jv/YndTDsZFnXOOFxbEBk7WGYHTj0LqR2W2GVx6TfcTixCKl/kbBpWGD
lrXXz6ei6d0ErB3P6pgEqpX7vT6RsOTq/830mGe+zacrOHVb0Y35/oSOXrezUHjDNFrZdAxkvd7Z
bF6engLiZHhfSylDTI8GAyIi8WAhBrmT0/hdm3UslNS4ECpX1KvC3khzo3BU98OkFQJtIUkxpxJv
xf7oVwwXQ+eVRl2IXnA1TX0h/MpVVOOUhLFmhoLpZTkAc/Cwhzr5D4X4jyIFXIidlporkF9cs42/
0E5BkSAd+g5M1AXyo84RcDG/Dw4RMcQO3gSsbZ92HOVuUlXtuADwvTkKCdjzQRBtHg8sG3bpKrLJ
gtT9kV976GTgSpb0W0iCKx7ohG0iJNQUHZrmctKB6W6oSF3l/32q5LWdUrg3+c6F0QkVQt+aQLQU
XDieuLbdbgZHxKPo4Yc1/7AqGX4FL5lMsh1pmNDOVUX+pg2+uF8s+sjRffCDh+Vc02CxweG3tR7K
OklZjIwLG3nVHoG3EgIVW6aAD+KzD8As7kpsKozOOYJCIa3nA2NOmm9TBgAhc4KqJHBk4i5Ee1lp
ke+t7nm7jwlqeitBIOqxYJQif0Pu/wDJf30dPqB6VblUTVE3x8c7GLVIXPeDxoGFwz1NdfOou27o
If8Y1XugM6H6AzlGiGAj4+dKfv6UAqWMcmrFWBIKl9OhhKXokraqj+dnCY7y0wGy8qv5+zawaEPV
GB9SKd+LdBdvKGCd21DqTC/nLeCAHoPagvuNwETwj6Xj0sNxenh2nncQJliJ+XsSeYOEQ/E5pfFi
x5WZgV3BqrHMMd6d41xdfLQNipoNHSlpXlsabCJtxyjTi0bD9Z1edHb75GkpKJga3LpJ0B6eRtge
XDb9+aEMzkm6U/6jCv7UAuntBGmkSUA1D5uy/7tynRWvmH/UoKC31AxPDs9i9p5fQ96wODx/eGMs
kkjLmVC1nQNaKaTGPJua5RtjiYK1E6X0ag2utO8uP+hjtLLpwRwee/HvQyo2EGy+BXXzJjar1YzI
eS0EObNaNbimq3+3DDk7M7g2aoZndMMkwBGCiAd+JsLmVDudyW4CamkPgQqjBzcntGQfHLS7Bd1X
HbWJKhNVxerdKyVKrF0mGFzOA5oRCpKAtzKrtAB1yW2qABWDnijD1HRZibLz1WCHJgSuVVIxWLt9
GN5ny/HeuDYkHKV2hUAyMo/IyLwYzSGg7TqBY0vyJKg2OzQLDZkCSxIW/OVoDEodCYt0nRfutiLg
E1xZJVBr+ZeqykkoAmBzJ1z6ohUASSEZxy/CEENsq31iiWT2ZfbFKSXw6Oyy5cOcRbg5Iw87qZKE
uxgxnlL6WMALakppkgjZ/wSFZiP+Wl3wRatoTBD9LN5FbAlgJHyb4aeprTU0tBzB7Chw+IFWJLtg
1yqhT7PZPnc8/CMqgYjEd5Qv3jqgTMP8fM24kqV7Cn8bpb/YXD7anOaJdGNgk0sf8EpIOiSqtgIW
bGmK+ZavcKNc/L9Hf1nOXEPpySW9Vsctw8Q56iMWGb2f4TW3vyttZpO9f9pvPlyAmDgidQgu2RQo
VPWRtC9/L0ne/5fpno4K/cw49namE8Sqjzz7QD4yXNC0CZ7Jt071HTUX5M2H5YQ47YOe39dWDfBr
wDwGcQsgAkK+HQ1DQlnIFjyHMFUlLuTdU+rULzu6php08Gd/5APKx9ROcdU5cSRQpwrZmY5uGgly
ze8CU/njYIo8MOcTyvCIi/vDARhtpar4JaCakElMSyAwRvVWU8rKkQDMZrzr3ssjKukfL9BcG1Gm
GaGKFfD6gqr0rSXCGp5PyrkVe+D7rdpXQdSX+ayLZ4fLTUDuOcyox7t1QUjVVDGSVM5AnYtEoUG0
PXhIua0cUxvhqa1F5uICKKdUSVjdXEI4PETzetkEuPD+2mDguHBAmC0vsrnw5fvhRHGnn2KHl17F
FglGXFyyVMycxhEZUA0x2jCumXzaGB426GzXFEAg3FMynihW60p7GZKJO9Ob0xvUjRGE7hGlInaY
NX3NCUXZJjRL9xmvgOHwAs37O0QFLHbCOdYqemM5KXqubOsJw7Nua1jAo5+8Y1a27zhvitokPBHt
ORS8Az2p2EN2R0qXDXywsR+PJTIqkB5C2GkJv0fepFCNvagleM2u0jHOeJLYkymaLKBWMA6QUs10
b4WMmzeClDVHQ4dw1sRBCpb6fYLV6d3MV2Vdrinpdw4Px5amrcvSY3mkGpH7bZXr3oisSyfWDS60
xE4STkxO+xaVlquLJ+273gPCRutfoHzy4Pr94Y7/fmwITbnUwnF8npXoHwLH1PRYe2/hGJLoQA18
DU+q6H2acKI+eV917WpVrDoFJSSGsVPtUYA5eHp+bOXO9Y/pqMHiL57VbraXCML2YtgJa9WWZNj0
XFmhLvkr7oleSEC/TDo0p0vQEbKLbUjp3CK0xK0LBLR5p1O4nMNBOEaqBIoLAKzl67IO8i2jrAPd
632iOcbp70Y8KCDfH6tHEZv6XOqnSJPgn7cbLU4cgZK1IolEPTfRzjf/p7oAnTFPBXb91N9O3PdF
U9aK1kuz59spANt9229ERMbhUo0UnJ5GmtI291Jdhn5+iHZr8CWTeUzyLWftt7/V8MX4o3uwpaKq
s6UcrimJxxZVaSnIvbrJRcLwlF2Ubhq0i/PWzV3eMW4j8fV3ainqmuevsQkk+ZRkRAyCVxHBoXy/
ptQJDahKkwu/DMg5L4rwQHo9cdgabNw9JsSUNa7W4QHFukPehMGg67IqJKkXZzrw3/HgCTu5nKdf
KNw9amkkyoFLHdisT9VBATkITxYdbhOQi0e4JsKWa9c95GN34nS23/U1+IFf0VkiuVQtnFMW5kWF
obI2n1CeQDtQ+pf91FvH1f+2A2yUz95ZdU59/DpaR7E/NgB+hl8/iNY8lacl8LIaV2CoL2L1/cSv
edgyrEC1SyY1qsXTNiVb29VRMGIFhssvXf62FBhN4CyBb1Ul3p9eZdh147GRSmTbT+mA4R5DJObL
Gl0e3LvA9GcLo6SAO5c1/1xCQhxRvgLna8JjCrJKB9EIs13XetzEZa6WhOSkZBpkqArEWT5spm4Z
K1tThL5EKroP3boFsC1YpP1poptD7pHx83Z8rxkWrWiOwtCTIV0YjrUq1yZhfOGa4rfRLb7yN9vy
cvjXHzbc0DhK1U3ozVs3K0ONznKPdOY5RxKPA+B5QbOHs/dExlhnxqAQN+rSuT1GF9/bbhCoc/pd
U3ug+oBo5xRa8Izdr+vmeyxoJfpWv/Xs55bEOHRNQ0XbMYthS7/s8ymdNKE4FaS6Z0s6cHb910Nt
pK/B5hHbsGBRJtlkZ+TewzvZBlkSgydVAUnw4horofuqy25uBTPpi3OgAiMcCNcaK2zaUbjfVloA
vhrAmRxOV8DHLbQSOYF79PtuH9t3qHD9r3ELktnNr6nouSXxeSSGdbFijSvtQiwa6ldzV2b2vF2/
Zi9OoqkHQGd68kOoKbkZa36flqAJJaWLxe2mRPxCGj0JaRds2TTEP7INTOezxjppVgBWhk699uf7
U4dS+g+KeD/MSICjUNvK+jjvIrG0GZPJ+T9mHs2leGWr4W8dO+SaDqE/xJvxmHPjlHqphs9mNkuz
MNM7xqH/y3PviRpSO/CklLl+IgqJJ6i4eBDxfQyUQWM0/+29CrNs93bGnhZg+5O1600fwa9Iu8qN
zHIyC+P9Xlcxw1XA9YVg3VJSO/0M0l7spZ/7SN8rRxdDDbva0z0BPyamtmyLRx/ZnBqwWBa7dwX3
8YmzX69lofMq+gsJl7cUATN61/pLeBFLbPA+quCqK2bAWlPBMmP2yflBKlXca08eHjBNgU0AXkKe
niXIavdk8Bm8r201tG6yDUEovSQUrLTWeb8GH2FhRUYIaJUq6UfEVw7Yg+badfey5INIVMw1rxOV
PxNLkFXownrbB946pIgd//9h57cAqHrES+U5lk6q7KbXMZNjuXkLOB7QtIvtsYmKG5Rw+FQ+HQid
vyGEF6ErD5s+/YqidV19LyLgMg9v1aGXFkIfQdET/6eKZhPr/3oCMtZbfOQ9/y4/mzKv3knpQyuA
WtgbxSvOPB2or33iIJi/ZSOheneAy22gdZ8h2POH0YN5yqq8kRZrMUSlxnM0hve43Fbj559shwdY
cs9ntojYHx4nces+QVyY96jMrz9TmOGWUUQWWJt4hyh2wswjwNU3PQD+D84WYRvhNZM6x0PK1Z8B
neEanARl2CwpZIcyROPJNrXK7vf0TSXuPWav+xCfqBYejP4HGO0oBidLviwQQUej4uoqyVeMqS6F
0uWZeVJFhkZcONAhFKXBS1w3No6fBE6FPcQRjepjY6cPw36kiOU2RhbobHIOdZlucSMc1fw15rTN
EARkagOaEQybvA6OqZGZVVuQc7YKmdzuTVRex1ekp/sdY7ru3dMVQVyOJK6VCtdeqhT9649gorek
vrtwfHZ9rGXjD4FYdApc8pL/yt9CSNnMt/8ItyoKOnHnxP06Jq/k24Ze+V1xDaH1TUkb+sHeD99H
4iWnSaA+hi/oQ0kJgay1ZiTwBrOQ3+ufECv1tsvZvZ0IPbH7ZfpcoKxcT8OGKYNmoqX+7KCoFKqj
F+MHmMyOpRhnULzn+GJjVYciNoR25Ci0mldI9gMWCzYTVj/UibqSyff1EM0zZLGU+gDr5eVO0XlG
af3rey2gK7FazRgbX2I7qJaRj+Aij2MFiQpPz9uv21N7drsfif8nOE2tYu62YQwGta5kFmM26hox
asNu1BPYv1gX4g3h1BFdb+2fiMDtPkcOO/YKfwBpnyy3p++D0hTtNu0EVokF4YniQofbKJl78VWR
2NPURF/6xNosHLqfcWKfuiNzr/acl+Sgw5qpXDOANKhT+Zdjri8JYymJRRmi/u6Ev6hUYKRHlINq
SECUfRPALtK5V7F/RH6z9frw7X30zYtUSgd/UlCHt/fRec29bjVME3o3fGfNCXoM04Ks2kUKP61N
b/yuPDEuTjlTqE6gix26RGc3xFAXRb0YS6Nf/R7z7trODwv4sZWk7XRtnqk2maH/4zLdOvL0EOZn
+d6cWEci3Xmp2w3UF6rNokyFQIddT9kiKsUa2ScMXW42S/3VzqBWWrK9WNVuLjdWAyfm2be1u+u7
/bakvfw88cxC6DHHUGYwpdeEqlG0heAw2bGA8diGzghu2NgGkVtBViVX2/D0xVQ3LV7i5Ji7df7e
cgn796Ag2+XsrJsTATur7u3JiJ40qfbLFkBoZhptEZrBKLa7ZXMALEIKXZYE0sVZNg5Rx+Sad0z+
UB18nnfcm2nhHETHz1j8Y+jPrMtp1HJrbgH3YCcyuOY55Q6r0JiHljHVDpa1Az/3IfvvA6UwBcwk
4C0xaePc7ZjB9exxe5iFu6HHANgkPA0WAbAOenhc5hqdBn2ucZmcWcZ+uhaeARpbwI8HHIIfG4r5
tDKaqspoj5dly0IgBcWPEAheBIIf9QaU8M5wzA+03klFynaRFbIdHqg+AjtBYK+KssbnPYMQetbY
rYcFyumG3rM0Ih8JXfRSdEPQyWv2J5joIYm2EvXdGc4JA3A2tUlAJLROyxop03vu6xd2ZHcHCK7J
VbVv6D8ywJKA7JoygUaVQGAqTEsgvdljCp2dYKMwLRaUxrlibgUCuQAVnZpNUk9x9UVrlsXXThUg
O/gDR5bB33xQ2+xq+eyM/WOGjX0uW6cKDyTmvUGz+MB+IstzsnxxmZKgeatb1bOZe/CyUsQU+/Nl
AwL82mVhjWjWFgyzwjABLrth0Lf9q3GSE7qythIa6prVa3qFMcOAmMzic76I2Eub+heK3ELuUsZ/
fsYbTZVhXJPgwt9Cxxd70holTBB0AqWAeqr1mK7CkyoJPiU08F3dVtFovZgV+UbwSGm3r/6lC9Vb
pnlZtC8aB6oG4HDfTVz2ep8oJz2TZKqxkzaUcyeheXBInGEuB5oHzAiRo0z2WIRecTCk3qcssUWy
EoNwsCBJsHpGamzM8At4J5Q9N2CKcvmAPhOiCbTtZC685SPP/A9W+dQcdof/B+f0ujdgKlDJkw0s
wqkIw3XAjMcSdSYilFZcyHy4lQVQxsay5gB4JvyYI4JqL9QKfqqFy56lZEY7RJ9UTjROmvgDYDlh
v8im9AKTBQq7e295ZkcRbMb5RXqaUjiD2BY5A5R6VB/sH4BPb6dIyluYZxA/suVy0p9NDGh+aN3Y
FpNLY5Y1V9HJEjD0Oih7LQwYH51Wn6N0ojrkHV2pV7IvXhq0Lz05zQQ76QLDrvHUVHsrig2OTRKy
E/zpdmLMDoA20Aqhp3PTwm5rQ7BAf7qReI36lEiYN6g7Vjm8/Mome4mjoXOBD9Ksn8V25uHjz0U7
lny+EJKohg4GpDLmIAI4qxZrDC7zUjQxyOcxdK8QrTOCg3EX1tPupMXBHLkwHK7UKkBn6sgLlH5c
EUtLv20Ka6xc9Hdckq4+nkztj9cwbvp1vcKhSlUeKeiUy+B0WZjz7N3qvhO4d3j1AqDn84VozTZW
r+BkKo5ArTyWkw00wxKbc50unTXtnRKeyBVYDhEd6VpM/aVFSFamqhL/yuM+5fcF5/1iMV/DTX/K
W2YbfN7+ouGtjog9oNab7mEfbz07avHMFL6J2vshokEPRMJdK4gp9ekUh7WGqxIAOBo1rBliD2yL
HbcTfW1w3sGzfTB/2QnRWKa9oSwkSHNpJgfPA9uMi5Xjf5OrMO6En8abfblgib1k1aB05B8gw+nr
NrK0zBaT15e5YyhAaXuqXWPSrSXvKpalJJn0zGYWGtFM/4U3WmA5uAk+8W3FBRlWI+vZR+u5/Bvj
XoFkdThkZk4bYsRZgXD3TDbGhLc9kWFE91NHKjzq49z/C/QejuXUg8LC4u4cRyCDXedwJp3FwmRE
MH8KJWxDse6cPpQPv/zZC38NvwQT3+t8J4DwtjaOHvlFCHI3L1cDb9LEkrj2zxKTaNTkRXUrUh4d
cbeS55M/Vt5uq69gu+t13ULutnXKDcB8V6VCU5QkxwdDt5dJwuawRMjcyI1D6DpwDC03INqMPEnC
EkxQ5rVNL+NJ9nRn9wePEqT2ugX2/EIGKso8CaoRprtrtrtfy0k4N5tGwlCx1r6euOwfF88pntiq
XOCXJQiNBdlbPRx8TMb9RjBv8Q+VuX1yqMVjYlInnQGafe+mlvGudaKFj+aZ9PVKFefQT34HYEqk
pUgyQUOQuIP4Tzlva1Dy1bml5/pM4blf1iO/e+BVNjTgujWqQI4yYCoNs5Z1EBhfvQ+vTEEPvRdC
iiK6ViAgzsLAfIVhE6Bk3wb9mGCm7oXjjIg86gT+VXTX721WVBYSNcIzQIoqBIh4/z/FmWxWxspu
YfYNUD1eEsAJp1x0YmjKVpva8Q7XKvAfFry7TyKAxXHfaeZlw1N9IqO60t3pHhPLy9zN7WO6TRui
fnDU1pTW/ZsRVKk6R3tO74MIY3cSIoGpNdiMevKlVFJcdcnbryXxU1sblJOW7DcHft8EA7mIOCdJ
GR3irM2ZDQqtVmZ1YUjVvP8vIuyFlhlmzuYffXy4+FpYJX7paGNJllwc7WJnJwVD2oV5luomlfO0
DPM/CM92epjZtBZxC3N05+sXP4aDld9iKAiH0Lc6UekRYB8wGGEEHspmbO2k1nvR4HJJlm/SllGI
K/nIE7HXxzXstvK2Bix8y/Tq/mQ7fMhnm8sdStx7FUcFskYHV/wJ4F5u0gWHKH6/lBA41EOLIiFZ
imJ3TReVLg1XYnmXiva74J+bQmUhmGDFipxTgvxNOCzmgU3CYAH6BPGa+gDHpelEDqRKbb7Icoxy
LPCWstGj1vFFtOwu+1WGV4TcInMY/xULnqSvN17go5ZdgHUcdoE9bMHx7LhQjGZzFRwbT45oQO0d
KHL+3CmFsKM9d9/uXMQ1dfSR4y4AyiB9YHs4X5Zgpd8DcDRjE6JBlcXP8TSNWb7TmIjawQY8tug9
x2ZAuFKzbsuNzBYZiWvoP1BHgiyYXgbul4nWVbKs9h1mhDpkoL8z2WKRV1U88STmz2nVHKI9V3/T
X1EgeTqNUrrUi5uwC6fV8VIfGwC/OXluIdlpF2MgIPD6FfqeyIxku2OPewBYzYQQTmsKJk6vvHD4
xjk72r9cZgCSv51iB0ypriyURS89YdPttNm+1oAcSsJ9YVM93975F5aAcLp+d2cUHrIqvAVipn9W
eTtu0mAjSIpQoH1g6AHgEfOis5A17XIQo6B8U2FqhhUeKTSS3RU61r+7Kj3WxgGKv+GysKFHM/YS
8dpOLmeUDxwMWTSmiTiEoDIqsS7Vx7QzSt3e0yP9p4zMyPoCfZiSPQSBBBDEhU1B/qLUdH66xyK4
slztf2Yx83cw+nfGtyOZiR0p0GelY/fr9xBBo+MsoNpleX4topWqpGsNri/TqttWKxrkPQP7u3fu
I1/lnaCY+2SqD6amuGPNAAYwsy3x59X5DoagKPJobqF0SQV4gzTwbBigCqFH7amzNLzfVBQEbuQK
orRLlgOKGEJqgz8NAhgWOyXKywsESUi7pa6k8sgFJ3eja2sauZWGRSskt+Uy+g4HpT218Nx9Heg0
iTKk/Wh+wr48k0xlczezZ2UAIIHOYyq/uE6wAn9BU3sPYfdmRDvZE7N1W3mRB8Vzhgnrt6NkiARa
iryfjIfrde8bBXK6lLF5IZlykuNpuDLCx2nyIlXIyYB4t8J+VXB7u216OsmGbAr+NcnQy3DU3kcI
PqdkvUO8TuxknrbJKf59mI+vhEtAdYb5yEPv4/sW+qAXhIFBLTYCqMoU9yRU5fNcG71SJl2zzIn9
ZI1wlt8OA9ajGYmlQGhrhqVAad/JeNxwRjFS/bX8TStSxatlUAmfhTIkTEV1LYTb7xXGN1B7tZCp
97jTyzmORYWdAOYvWUiAbhR1akIUyeJifgSSYjv3kqXWGRABh8Zqso+OnoUEd3Msbjt+tVvO5wjq
4VJoZxH9u4Zxxz/+x69PIwOXOda1ccLHeSqDz9s6ZFxGHOXZnLtqZX9QALsHA3JngNcZxPq6ZSje
7QRR8KgybHzg4+5YnmtLeU6eEww9WqikUTjjJGLE2yf5guCpWK35pCWtlt6G5f0xJVuVLaqf+GEt
t325q3baq4Rs5AqHXDgwNysb2pzlvp8XBE651TgsEVPCG1x9cS6T2JuZQmlT0p92+Vskzsm4KXer
hFKRES66rzLzOcNXj5ucFLOFcW683C9Hvw6psMeST4NTlx9iTHtSAVTHhwN5wj3ixnzZEIknu+Gn
fGRznxI490CwbEE7RwztUtwsbxHYe1e9hxGsPldRfpJkoCgmZnYLEmI2eAmcRcKJMc3EBhzT4urj
XMtQ/Q+oQJRO9JXKVyvw0sBcPFeE7P77IsnuPrikhPEOtx+E+MbwMhlahqOW9BLD/jDY1B5BS5Ta
g/6iGinFvBi4vVPhpW2tRWAJJe+p/8LwcZOYWnaN8DEMIWLxlA1FtAMpap1vx2OOJTWTfv6TzFBh
1y2PlDH6cxHF/kERgy35TOg9g/B9dEHV5zYB9xIUCGM8COEQv/FqvhC87hn4S1+JHNutAirLk7KM
yEPNRbim4I0mwzdKfml/OOqg7DMMFZVJ10w8hhp9Wb+zaFRpuiT72+XPQGTcw3Q9xBNO/DU+xMCN
e7OxdBNVYG2D0BZitDjU7nfK3EkYl0KWlM/tLKKUNSDuuS10qDuHFOfPgmwPz97jl2TVLUp5VbPK
s7WgibDqF1uQ7Ryuu9Q0SbntxzOmm+8DP0BR7kxzaaO9q8EBNtgq4mqoNfKIGn4ams+kXlKSO6vR
bQuegEjHc7q5dq7rvvFhfdjmFf3XIxn///zXdPLgCQer7VDud7PJtQ1OXrT23xsbE6nayEt3FrDP
YhDd20ox8/51MFX7L98LCkDTljobPxOjBuULSdq75j6aCXeBfD02QjIe8Li8mkZw8gdw6yUQXr1a
tY11eUrPVthZ1NenGxXi6ZKyjCMUdkhXs9CDOxFtvAZYvSevoiYVKvCQxNRC2KuOJaFAIssz5rAs
dBLmKeHuK8j+iI+OA5MvOc+G3r2FtAdi5IPDWbBn0EjEVqzSBKU3sa+QH6QJUvDZf6khnPwXRRB3
pSJFSF5rzz854PUzAoFzfEBJ9QCM0OZFz0Vqbfpk9u4Jqak+f73Rq4xpxRcozeDy3GFY3ra5lXyF
d3inlvpCsI0rl5LREJX52jWuctXV6Lya08eeWEayqZe9RZeZ8Gmb70l4Cl5NIF4Fq3aLTl3o4NVA
0kIXrJk6frKg28j4LqsReeCahHIfn7r7QFhonSlOSTCx6cAWW16jjqGy+PcsgmR+RF+wfPqchH74
wT/Ja6X1+NXzQ4cyvZPGqH+iY/VHXFZw8WkIT5Bk+LjsFM8sFVfpWWyjM9WK98hNUo8+gNVuVBZF
+fk5rUuVJwckZLgINZ5xajXaR1cSwMtyB28VBMmvOM1UQbao5dss5Q6nv3BUH4l0QRvIYVfnGeA3
X3r0s9hih17Jy0hvCP3iJuADR28OWVA+eSk3mERP6ix16jkDnf33LAbJVljn+P5K5paX7oGEXZbA
xmAAD6h6zINPdnf4hS09iVdnO8MX8FPBHY3iDb9QBBDLADbiMcTTWknZT5MQbbTxxxd3keqclcQh
c+jsKJY6yfmL0FlUH2Zo6E+o1PA+yl1THd4S1izpa8AE8OOa7Gth53jS4J4OgIpIRvb1vXF5CSfQ
VgzTvnfujcwfA6e7eJH0fMVJH6AiD/d6DOHO6XIkRV6XRhkM/j4SzxDx2elr99Lysyx/xpITptzv
MA0K/D42OPD339WRA3OycBPrJ2ztMs3HQFude3iHg7z166e7ZYK0tfqd8OnG05flLIKztyTZS6Jt
96VVNfeQrlXjl/Bj6nBa5i40dxNgqs3s+ESzEWMmp4J16QI42+43UOAHfBgETBcYWj/tshpsYkdU
hhJVQBCR8jAlAwXHynLFLjYVhrfds11CtJLJUBy9QCkqhyDdCM7pSoD5s7YNIRlPC/lA4YsskrIk
wTkfAAKkbgM/VRKlNsIHBeGlJ6eNvKocl0syQZaC/+SKV66eCV9gGEiXnBZbQOl7XlWHrXArN0K9
+qbOOn9/09N40oDa3E7Qia0+sVaxpWLQyWZN9xK8/tnMhz536WFUsy6BRcY2hIDix4moG4x+CWsn
J8BAWmBaxxd1w4RBVv7EUSYlZy9aiA8UaSyLd72dNVYy3GV1/nGNbA7RZIQvYV6wRiXe31q+y2MV
XGC6pggv9Hp5NKQCK0oBogQnJYgQYZiMf8XBR+DpzlCPrdakSKD8P+JrGkzavjjnveQHpNWxOfGk
+GON/niZBW4qbvQ0SR3hMfBW20/YcDN5Fu9AYJclyP4+Ikh1n8uAV8QiTqEoQQIW8Uzgb6XZssYB
emEQaNM0k2FP3mE5PaZsc20IbiJf/T3kts38rZ3yEJDK0iNlyv8zG3z5ALMhxGWcja0tBeNxNhas
pzdVNNGGqeGovGT8mAo6cOJY2imLgj5/bLgkBCNqzssXJS4awLHOMHhmO7DfDIqmgrfKXeLpOmAP
LWqIRWKrVJIMtpXr7oEq6vV46Q3uYCxFpPJgndBp1PZiKy198vB8WEOjvQFaXTkX/I7O9GfdwI9T
fL7MkEuWJoN0VtwGCWky3Mt6bnu2LQy0R3tMEN2rkR/EIVXH52jCT728wqOKXJBKharSbWl8GrAG
mnN2PZ668MfdmQct0AkGLpQyEA7dlaFMD+NNZGaRwZ8JgU0zxIgsiSNuKcyzmIboz8cbPZYxoADn
E6l4BwggfaXtgn+gKKug6xpmMSnQwXn0iyz8EksWE5uLettnnDcR5xowEU4AnWHCxdXnjUINB1QK
lyuZVqBFWAt1l6NJY0gf9rrwb675vphBU45Td/GkOROQ8MlKY+iug8gZb/NpPanbd92UXLDSgPy/
rup5frUcqT6psLlz3Vvsmhzx6lbU3S0QpzSL4Zh9jiURwPX/xr4dKi+E7YG3UWkeXjO4mN+zHwFh
JZwIYVQh1huDobVIY+amJyajQfkyDUYb9zHrSiy3fVNSDsLMQ2wPh2MlWfkaD92mb++HYXAuXZFf
ld9TRQIQefSicLqCOoU/LU6HDNSCpvCOL3jSpcerOrRRH7tiIHfxw0CSZZ+SGyEh6XoBftxpSzuj
WyEkYy2bTWfJxsosNLYoP3ukIo5A7DK7UfXJRBO7FotffIhumP31DYvw64KKfVRht76xU22eZkzw
vpKvBAiJdmTEKJRvIghf/Fzp0H1xIOqPEGw+KD/Ggw5lpbqmOCxqL6YzLQYMmip7/yZlaVXOs2o8
gZZLBio2hgtR9wFvrr4zBjHhdtFof/Xw1tjvL9BoG9vAMlBlyA1g33VbKuWEel3ZgQWUvCB0I72d
SV6mbjDihAAXSWdlQc4kJwTgWRgwOGMPKhK/fUcLEPV9nV389fsbcMNIkMhf/eQGhSj9HNK1piHl
pbpuS02rI92apBI28HXoSi1g4Y6RbuJSVkgdB2EyR/Omdm+E+ceuCwP0j2psj5RJlzeT5IYyQ37C
SdyA826jXRrubCscVhJi6O55zgHSd1Df93gNJeS3WtzyzdvnddJ6T1Quekqvdyy9CiJB+GK1kMtA
utlfqjbxL3aZoF3+beESQNfeAxFKP2ivCKGc8kl95JuyK+rKzqHlgbkSGrdm5dCF5t2LNvTds5+r
ZgalrGPzPNIZfmggzVFvS3InRXwxcyxSjR3gB9EeXsM1VEl1VQNt+6dAdSu8RbYdegc9IAUrFgTZ
Lk4Myuo3oG0cIZIbk335l1DPPJ8Xrs5fhWau6V5Gm8G1d1JewEmfx2m6669lrkUDA4Fc+5qJ16ig
pv33rE0trK+Pzd7YeN0CO/64gAXBYsEKk+Da+gqkkKspaVI7heF013PDYye0cYZXFHjzS00o4DWd
MnAigGQGFR1liIoDFMtviPlduyB7YekziVMWMQzuINdBI2J+orJaBbPmuZzF3d9iQXR9ds1atB5K
dVqN140/nQaCj31WW/YJU4fL20uEUS4V8fu7mphC/Il/XXlndtrwaJCNIBLxA5+F/yoX7A5E2CFr
LVpNVGRy+UG7IjQgo3Waciyt43dMhh9666pZ/50wSUYc2SxLzj0HYXa6YNEqzf3dAV3PCXb5DOZd
d6ZFoSH2vFCKmkLyCMmfMiSh8RI+1i9PWPeo348hhR9BFfY7NAHuEj67IU3re6EK7pQpLGYnByaD
m1dJB+heEW0FYwOoEzntTCeIF/f3zk2HKXYE2sNqTHSgi3kmFWKLFRkJYBoW4otKsK+kBUlKGQVs
NprOVT5wWraJl8sT5NHZSrkd+8vs6Gn4vwBCSxqzchnEzmcUC1Ld72sq2N8IK8yiSqv8B+NKVwqx
0XmQsZagjY5nUbyGtdYSwDOrqA4fsJILj/7DdI5akOC4tGCYy0YlfUewHbrA5GVYvldNxS7tArpd
99/FON69jLHVfexVQB98aA9IM76qNpRIz0r+88WGez4gDyRsvaB8EZuLOSsXhDrS1Y0d7gNl0Yxq
VHsetFyfLNT5f1cJ+N9gEN8c+14MlAkzmgAISSalrNlpucz80yiw4l2NNdLfMAkFTVl8yfAxLWVA
nTxZCHMvSUA7ZMdC0elUGNi6xO9Ax8UcO239aVJPd1NmW0GYnWnZg/iLP//n6qHJ9sNPA9c5zZJj
vbA1ExjyJBDtorYkTYVy9UctleaVOPNW10nPXTUSthR1IJUERGiFUpZmK6Q4UV3/YWTIqS6yKja8
AIYTSXUs+HqtLzMheIfoCGcpxdSUYUjY9NJ6ZrAVWRB7I5xAfwsypHLDqyjyrFoT9aRSLaLJkarP
MDNl3yeoUI5JT8m9ox82S6fF+DuALq/pI8sV31AbJktRXcX0bvUAt69xSOjvVD08gleM2y8uJMjA
kTtNkwJgFZZtDZtdiqLAtosoC3T4JIsQLmGioy/LImlQl2Z0MMaJSOtCOi7tD8E6eOexvy5J1MRa
r+rj05wJ6wuQdzp33dJjCK2GeVCiFxjg0T2lUHp7ynN1tyyFCwQ/dfmhF0H6v6rT/QIDDVeBcO9w
BNXDiJEWziuwXie8cDwyTqvwNHmXG9F5dYDbQwj70uuSg9G+v73YK71tTmqP8ALXpX3EVzlw+3uB
I2K9whdH3QzDH81s/P9iKIDa1/GWZiOXMyNG3hrhBsxhQT26Wi8UupECkSajirAdOnqpMo6+ERoc
76KPO7yZx859nAAVyV2w5v8lNpEeY49xYvvn7z6SenDZl/ufp+u8gzLeIIztnKIJDFDtNooydYTt
k7CtBkGJXqc4ed+hgo22OCyBFll2fS+VBl4+Wb2Mp+FxF8lDne+S9l2afAmmADvyrxk/G5WqNVmb
+/dwelLv7jRBEBzlosNdD3BaeLPQqtMsXm2O2ZzrZHWlGDmK4HDIt7xXZuPmyj0Inl9OiGIGPtey
+qxe+GRdCsTtrs84rStGZRAvtaqbRIesNc98Bv0yVa6GxEnTsxNUcGo44LyZhhT5A23FuUCK1AD+
rKXj9EieyNjF1h4gAmwu7eKKTccH3Ir2+9oSGkT12NrJUzUiY7+K9na3YzMIq1wXNx6sC17BjKPh
khRCAeSWONsrWTqRr87wmVaNog6I6WGPXC3Q4+2Sl/anNvJFE04g2dr7PeyLvqUAuC1VO1plVeS3
VDWJWjBTXDV+74lr5cCUk2ogB7OPWOzKfbI2BrAcbRcCNXiNGgt7vC3CheCEDZrQ67TFetTX7zdG
EKwdzfNuB7xpu70O4gaiEhtq3yrNMjxI4nuKbyGrFjA1+ZeITKgYUBD+xbCCRC+afnarjxrdMhZN
+455vlFIwOeEhRe2YimegaKUTrP30xyJ0gV6BiFrRSBJ+2ZYFgS6nLb1siGHY3TmYRv3OBCoPf5S
9FSoeEKzMtPGy/r18x3XuSKez01NBTAQPDTrHjH9ZEYfmtp0aql6CStcZGlk5aMRE/18AQJiLBli
qj0iDNCWIOge+gQ5m4DCG1Ik79Xd9K8xolYFNhM7LP94aJw9tHLpGKvPfDTYAsyX1Fz53M6QoRxM
UGsBxtTFSy3OVmsei2eDU6lgaQ6Qb6SiiDfCkKwB7XzW+zdRUs5naLtUqPJ0rGmVju9NqL9Av5hy
2OhS3c+uOyRPwQ1MUx+0/rumkSAxEXldG9drQQqhZ7R+BKZZCn1qhDfmvwhEvcYRm6bgjs/pOkkm
3jI0DnYmuj3QO9jqARTvpr40MpzGhJ/co+neo3UumQ2BplZf7YwoTBMzRNPCANeIW9UNUOn8nW5H
gNraAY3Jd2Qb5CgdrlujZSyd4hpcYJXNVbTFqUIgTU1C+ig9uIHyo8RTbNhH3Mx9fjWofM42ucZM
TCfF67siPR163HBh/47U4i5K9zrFOEGLl1spJ9uqjWUZyrYtNnjA+fAB6eTsRI+kYd4QwmG4hFGV
u4wKxo/IDxyX0Rmvgl0xiR62z6J6a977uau6Y8+QFuNjnsXvOYHUgaw70Ich4Rn5d2CMFa1JTM+A
dgq0IbzxvRMaTNYdufqV2NfJhLZbx//fTM19YTQofLCv3aGsAAI31JnnQGHkvP0m1Xp4kVhE/k6h
v0C8lNnATX8nql2FxhWNRIgd3vlo+6d70+jt8l5qKXtJMfz0GcXJRiaNhE7ZFn0D3PBA65y3EBQb
7yGAhSeEmETuB5XuZlBWfg10s6NdY+52REv3fUhuOdd2dK1JPuP9ly/N/BqvKFma01dtzWjbKhqw
9PW6tlRzgIfZXobiDlbJvh2R26bywledqHhXguvNW5WC+Dos5THgDVfgFlZVgpTuAz2VnhQEZfDi
2m9e2WKHg0wNkVMY+u4h5S0hhmPcSKkPjV5kesOxNM93cSHKi4ENMrMz2/vCvzLUmvs38Ey7dh/a
zCf1fwkHEhe6sUUwa4afxOB6zQBN98Uype22AvqLX/nWmhjxnbdTEJPo2uloxZwzsxWzhgJvPFh8
PoreSuiDRUuTaasup2SMkmf2lXqveKIIH7+y02auUzG8Vdmsd1qPxjfim8mWYK3tf/VfwRlpok+m
ynby1Bnbsjkkml1BKNSOmn66/tnxmqYJ3SWmE9K6s3nx1egL/BKXuaJGsffQybntSjPVnRidgm3C
79phIPSB1rBIggmcc0ub+9BSL6n5qT3xDbzElSfqav8ik1d9pKW0viKuCWnurXzGMC64rkMGxcF1
RsQR2MFGj88SAGOXnaNeyY2X+8GAbVtIzWqOs0LiD5QjPTkMPioCOb+hbmQszbMGPyb0+F//thga
+ymog7nBiIR3fbcgTmC4tp1SXtYaPa/fOH+GF3G0WzCTqchmleoEMp5CXuIupKS2g44hOC7YGL0l
AEgyJiknxU3Z9w1STBRVI9nca4pfWPMHzad3l6XWTytg3cP0xlaPXE1lue5G99rql4w4OWOskrow
FPhvtvbuHxuVNbzZybkdk20P5NqJm0Zb9uwjRHcwgeN8nntWREjRNPgj3ROr4iyJq3D9UlOaP6QF
p3DCkEsROY48DAy9f5JURjSDlV+K4I0TOdWbyIZ5zhUeOzCxX5Mq7EH2FjQA95ZSVqB7W2snXnkz
lrxAJi+L6O73EaYfCOZr4V278d6ZAO9QkgVsHeLHGSuIhd1azGrD0EFDZnnsZtasuUb7oodCzVWu
gae7cAKMt1eT17IwgHCAD6t2THIB6ba0cqPIS0KSs6VVL4yM5OKxv9nGvOdbKlyg4dsnYhaeeraz
gqxByj1qp4Ly/QbRKoxWp3QtKXPinNVdLZMDpuW1QtUKPMrNcM/eNMQp7TnIXUSxR8Rq/mZdblIY
XyzP/05kxuZUClsNclfsHeKvMqCvSfM0pVczOizUSBe0Vp2tSLxRL5VA4yZQOP1kJvxIUMICO7tk
MzclDf6ltKPFyYWDGiEXgVLygNAE1QiGRGLYkJYu9XdAlrpvxqIfqECswVyVMit2TpE6MFFl14Sh
iyE72BxL3S7mxrf52u17T2jxiwDKHKsVkANiVqQ7+h/NQbhoClGSQy9B6klZqfjmNp4agCAzYNvX
aHIGcy1gvb7vVnjFS74+EwckfgvlyOrGvAnJL9VSBnLpVtAytEkO/g+MBV0UffjQZX22RvGv6xT0
lv6FtPiEusFEl2z7IBVYFn374cLGFv+VgxlSxEK6sS+uEmeeLEsMegqSZpgfNZghemk5VdLDkmT2
eI176RxSBtZdoh6iuheyRG8QbEgK5wacrVmKN2L+XUOj4idR0JhgAnBSJEhlMf9+t8hwv5BiP7kW
O4WTUZcyq2Di+ahxfsJ+D+zurfmWU0wQzYaAFysrUYMz2xmGooGKZt9TKP/6Qkv7WYvl7A1DsXZ1
Fh4Kmy6CZYZ5pvYrLehEvXY0Vw3HSqy7uR8qXDWX9ws9G/LdLzVAa4FguhEyTlgS+etnQsqsGl0s
OqI+ytKp1M8sf6OtkDzxKKieNkhRu1xxEMNHLvS2kdmy2vJgIrEpGeK8msAtVhpeX0VUDsKMfb0A
Bs3k+mhrehOVAu1cAbfWyfRcycP14Gz3IfAdFDOHYV13yQlubAk5RTD1oTPc2gTKYaIczXmsQHwd
ueH/HrT+3JFaotzgxI/yyVvOiaBlzi7Sj7WNFWM79i8hehD1fruVdj+BRzNjUsGwDgJ/7SOi4+Hy
l7tqXit6mS0GjWdt473U7Ln+TTe0sa1GU/H5Iaydrv6Flk3uL1/NSPIJiU3iOffrt7dDwGmC+F43
I1XcJZZsVxGq7qO54hkTDEDkyq1hMUxqOc8hpPAH4HB27wI8P4QWX6z0f1UfYda2lTpNWhs5hbgv
rA7D0oqI2bCUXyyVH7/IqGbYyRpI0gko8gmwAb3sDlY3ewn5DBhqUFqS0fN4Yytsk+VKGQiGnegQ
1GXQCt1fgy7pwe/WqJ2Ym77iE+A42U5eevWdzvPP/0YRIGrGs5bXe2e7FrVWL7hbdbFkA8lkFRb+
AnfFAe0kvlhqGUfidwlmk7yV0H74C7PoGaFHbOw2u4AratypEszXN3rI9zBPXmnRgmW+m5KFGxhP
jG+DQ6Zp5vzCDuGL+HM6WSM9fesiRik1TkbR6Lse+j+Iuof+UX59yBQ2yTeIvOEN5XKP7YOiagtq
F2chOE49rHGUBj9bTDjt27o+Rrjiei7n/YeegWrs28bhTgJFLO0OBSzmGrYFUPFDpQtD6T4dn9tx
NyFBWuR8VA4+oUZ6V5Y0TNinBMBWVsOAIXyboqkaECr41n6AzDQGGke31zVc3a6nhPbmcWHT+ZzZ
2NE8iBC9tF/eYCwXCwBE13WTK1GoiPylEaatNu88+sbfl8TydDHgiTWZ9+PUiByQzyJNxiqEydkF
kGjTlofdUqvMrxh2+DEQe6pJJlbUI3iYUyhnZugI54VqZrRtmYVYexO1Vhs/clEPtHhlDEZurjTg
WJpSQT5pQYIQ1p11vZHcA+r0f6RdXtiad3cJwR1BIBXr4Nm+OKAtVgaf158KXTjIO+QPUyr6YnSJ
q/4q6DuWgq/DChXLih3WADdOScKwqWgoFB3p98agP1uMi3IzUT7PLcL/+Sp04bLnIC30IoSR/8op
L3KnhGcG6erPxkPcoHaJR6wSppmXy/G/uEzxYIv7lq3df0b0Ro/uLQ2b+L8aRnJ+4Zt/7c9L1E+S
KRPS/RcWj2+3oW6dz29IXEVvGQnOk3mrTcXcjfSvzHA1mQQ+kCmpmVje4/jjVdxOLX5dnNW5BZBO
f2qRjleBFXaMZa7gHCwBjFmGgJM0+b9cE39zKRIPlnQX/R6nlmCr6TgSC6VZY2/dr3WAzfWQKEm6
uodaVD1Wum7j5i2ZctYaCF+71INZmQmwz7wTHSuZFYvw4ioIBh+/d63qDDpS31eOG4Tj40rNzuR+
HmqZu6yFLCI/ijdcPevqacwJExck38Enz7Y18fuJWfFLxNzqOwi+HroIq0DC5DH3hkfDjzjDOowI
M9VPS0JGHCvv6YNnCTU9QjESvsj4M9kgcnmJibtVr2yCnnlOZ2VYQyJEY5G1hwqtjbfz8PgtCVTY
hCw0tIiY5ihTvKWlqozAwMzvdrW0S8ptVfif4MclCsSCsrYHPBv2V8i/g0zTjNcjZQDO9GYQq9x2
kNbW9kIPaYRscdcYel7pIx6ccFhhpXSiPpPyCEmRKflhZBFaI/ThtnHAQSc+NqtWepTo0jrCtK7q
q1f7IbqZtpy5h8ncoF/ZtDtKkWDlZsjZxeS3bX+cUCoDPSBPJbslhrawfvaSZda9E91iddfD+Nt8
GcK6xxvCV7iAhImFhmwUuBNGBjB3l/sGqoRGIn32ZLb3WBe/2Q+tk35Y+3nlIvn6qSnldZ03xZ5B
pjRg7VhIxbG3UxQ+ZXr83sNRhzswyHtkUtLYttDehMx+tR/e3o3CKcwooiPRno1Mo68mKgv3rpWg
JbcK1S1Zpw2PENkID3UDYQHgkSFKkCb6P51IWRJFjKwHLv9if3bsyu3VudSnfWiYNecILLsqtqmt
Du6FfOVXtT6dBUUkPCUi/yRPWYt6HwRi4YevzMFlVrKkYZrFKGjCqZ1vIYtzcUg7ExJ7pX2fmiFh
RMoMZEzHpvTYE7td18JHRiQhTQSzy5fAWDgYuLai6FwVFYdg6MVLEKDO4EvmTvwwjdRu0aqsrq7/
LVT61F8l2VpL14PoSRgKFN8tdATZkG1n35umQ7xKK4Vp7EKSQGKO8N+aeh5iZf1z4ELoMnnVb8LQ
w1CdxxrsbjEZ9daOjdHyjpRA4RL/H7d6vGmbrbDIGpIwLCwUiuJj03S3CpnHTxaL8z0SXZ0WWmmu
UloQoQ3hFSe7tvvRMrsuX4yjRLVFEzAiQgksPn9xVmXFPLqojrSYOjXtxAwPB+hATsaCYl8Uz4PJ
SgjQx5M9vQD2OtO+zDYDIwgFxYmLmozeZKcUEgfPPXb5PGg8pP06hGTq35SORV3bVyyELELSKnFJ
u1jAtyFc+3ORrqdR78BZXeX4hEeFreBhaFyyo8z+/PqdwIdKJNHmMQ4GyhEiX2/Iu76JuRqCnpWi
3kb+9KqeeXyflxoeb72ML1m8WEULXFsXKfmKQO8Fe6s/f3IYsLNyD22mmnDo+DbG5k6T1oqsCSEP
cKi0FWioWz/foAkvfrmzQk+41XGPJZCaRoJLxmPR1Dg7i7uKO5YoKGtz9BZOBmK9AAdZv4J/1ZmA
2jiCfN54ZU4ij075MQw2kBQJ0KvcBAwEw6epxEMEha1a4W0wgKRrOnVVGER8EM/+RAtJidM/ysvL
yxvfU12qATrCKJUCTNUUtpbRd9LYzsDqRI9GIb/v3W5caQGDI/mvZ6zGZPizPdVvxibVlcY1jkDv
EQeHsKkAbuZOFNB3cT/VmrCWywTPvThuY5TQ8f+VVBBhpz7aBIYvex1eEde/B1dySsfOqvcBeADb
3XV9pipsZRcuo+pyIR0XBzewhX6R1qIzgsCNJffRWSrb8pXkGRm0681eqR5d4bw1VyYUJ/WChCAV
uXQKToFyaUVLriT3uY1qhowKmLcal9pExv4uhr6v/G7lvwzDey0hFTpUoSz8YKi93LvjSjxhadQH
TsKTEpb1lHw8ZM7tIjPGH4Z2dr5VW4y/1x4J3uwgWyZwRactc5bcnNwsZxEONfJuFZU6N/fUDiAB
yJ/pJ/NBWkJNxMeiRxLRLbuUWBlXgQ9OjMdNKtpGyGW2fBxgKhUBcZAMhPqqBkbbJq/08ldxnfW/
p8gtu/ro+IRi/EsEGwdHQVJvHQBX6ZAwucWE24hKHaREijfzHnB12WaizvxPzzrUIrDIoDDxxhj2
QXpWIrbjyQExPTpSY0OZYmn+kG/FL2fFYaBsVTGv4HOocbwIehQd89OduomQ7UkUNB5ZiWH834p/
3wRBmZCFl4UwAKR5/yvJt5MMAeO+/4nOPY/ODGzgI7gVdX0lOJl40icQSxK+Sima6jgvy8e/BFpQ
s0gznySZVfEjYXKFr8xXcZvqx+tcVDlQMx42WLgB0IoFdxXQ/GGeBkljQEAsIuyVVBzThNSv7J/M
52IMoqntHm6FO6WANq5qlLhLswDXwDeeir9wPtiC/ciYgtemvJ+P7W6IPQKZ6zKcWTuMyKNIgkXw
z3GAHYGGizNKRwvgP3Czalb3/pLE9yHWEe6bU2l2243nn5ad6RTFDoWjtwAFJc1FFHELCWuMErsY
mYEsIKURugX9O4PbbxbiwNSZY7QjReuFZ2bAEJtRN23H/AEOoqp5+fglbCI5C8Q08JJaRn+FwjUA
2hVIQhf7KrojWhqBYAcygYwGbrE0N86vyTw3GkOCco9PaDCccm1Q4vfGBAt2BOqp2pvSoNtjzPQH
Jfm5BxBBAGhzfMo0kYPFU0J+j1IickjpeT8QGN9yaPJFg8reHGR+lsW/khKLhT1Ss0HJ0f89/Uf1
VhKVNGTL45MIh9qPUggvVF54JeqS5NSIxRh+Mi716noIPen/9Foe1IodggErUoTL4W5ln4thJ56f
6W/0vP3ITlq0gqnzwFEsvjUV3m0Im6Bhk8hF5ubO3ArTC5c5TFGBgLCrIcb+tZUPgusX+oUGPfpP
sb5/A11Doyz06SFUfEFA9lu3VxtrH45aFY2Z8KxSJOTaFSPRIG/qqHH3UTLvFSRLDBgeA/ztlAGc
x5PYta1Bi4TZGuOF5GUVmuvIoLmW3UxyNTKC6i1BIy9P4+hQdwvsT6GnaHQrA9KDx6WbfsVk6niA
oqngpQ7TUm3PCKElejYPclgm4JihymLslYVU9tmGPZ9tiJCGPQZUlBYMb2VW0eZm/dj9px2LIZfX
2s33p2U0br8iAImCKdtn/gw9F4zs14qAVTCv2sEon+vLWh7Ooywiu1y1l4w+tMVtv2HdxgNhNBQE
GTs2YBnX6R1U9BDnxWi9YaL5DZMmbTVUS0l2FC+fjcy4sBIM3LBe8Bw/vgYyb+e/VDGJyYifKYlV
3pGCO64Q4dQHBFELMaVEs+w7OJ2Hfx3C+or63ZQq1EGurCEDTYwOrmatEw9B1jBauxvVdMVvORC2
G+tjokAvJSdkqU5iGstfPR2EGF1FDSpz9WvmSzVB/LydVDQFiMN3N4LxZ9hzXsdKOLJactrAfJrv
+wwZvfPdmD/OPKYLbqjCXP0OGX4KjZ1mVgrUFmrFoKSfMNpXMIHVGq5axYk5zImSj9OyiQVYb42/
FvdFkUVsn3EnV9gIHxuwqKqjg2QIFKPhZ9x+iLUfqYoYDJfoymfatfDvWXy2axNez8bt/pJsrKaZ
t2Symgf9A5Z4DZh5dCcD+uQVIQ0Op+sjuPkIE2gjLQ02Yb4jGFgTYVUMW8OMDQwrNTn4ZV807aSs
/OpJ9CFHEEMtnF74bmVgRFWyDgnZzFEFh97sj1GBw7sQBKDJmZs8uino5jd0sR88x5Gcf/FlEaLn
K1egNBFYS1U6qXKWDiw/fLbEEe772jENv/+x2NhedGnB8mYcGiJ7T76q5JCq7P2yajLyAe4G2G+l
+5BTY8Fed4MZqRsphJfQAGenEbR8herL0vkQLMlAgr0bxY10kNNLNEYeh7IDIa0R61l7oA6TZNCs
0Al/mQOIk6n6ecOV5e6H+4qUmrYjCiryJPfELFP6SY++jSZJejXXbIQH74/5cdYyBFXW8ZX/8yml
e1QJjVcCo/CiD6zBijIuG8c79deg1icONU2nht9ZrwfC/qLlT1hgt0eFO/8+kbMQW8iCwaxhGdLH
gzEGwFZMoYqoOmhmlNnP/OWLVlOem9+Bmp9iwUdHmxBi7IBDXwxilALlBOhcbKibmjQbL1dnfKUK
uTwTrAPt7157Eqxb0fLBAL1G9LyB0onPQOZo4RxyFN3hokmRjz4BCHuSITljsmkqXVjcRIJWItbs
dItU2n+WJABQ4tLBB3ASMATcKDczjLUdgToVnZAsl3xoG50byFyqW30N1moCkJXXLKOJjFWxQSZ4
TzQQsJqrF8+M9OiCr53VvAyfCXRXy3qt2cFyJM4qehLdBQoovDqSKPFQeqP56y1c/Oq4kb/rA3wv
DUjHpZ/bg+KwkjFYmuXNDC7sw6e0b+S5ySsVsBWipMsPXHRJrp1eNXT1+GsFE9R1WWFoSjyKwgPR
gsqG3GLOFgJZyu4Zih0ed59C20pAcaY++NwLSBAehSrK/VBw2EzyI8rM+XFS1dlFUKBWasxVSpwu
griXhiYVipnqL+3qh0iuBM1ccyZM5T0A3r5QiqF3eb2zWCQUErBhOJnOo+FFhkEJY5m2khqYXe40
sBJ9w5GRr3frbUY822SVMa2X7TmHQmeth6RZsehkk3aBAYVrNL1Oxgcs1N6UYQeuN6Lvh4eEskLb
VQBnj5qgN1uYz1+hqu5o3URV3ugItNftkeS6Q62xetSyz1kQ3VLVtVcwDiUkoOWXvIbSaoyagk2h
qQAlp1FMtDMFwlUy010q1lkPHpgEWa8PhZ/sSnphsqyCQ3sRCh+NJ/hEnoDIg77wXvBvrQbxVIOP
jojiqB1OJRKTfDcemBT8neT3ZTzRLcS+kj/uzMlMWkCxJdf6FE6X0vN+es02hR/kKRO8jrbVWPc7
UhO6ZdxP5fq2FyZWXlW/RVZpj49WsMdH8AkCDMUUCqCgQyfpKw/ErQhyMg3gKlZIjW2+akzooItO
ONW1611GWLgZcuytqw+wAsmYmHx54w0nrFTOH5J1Ru+3sOVEljUOENEEAtFDkzNlVGytzd3YZ1tc
3Mr998Ptumg15QmJnCS02SYVPA/q0pCAGOMnVRPPAso4K178BkpkverUPAQJsRc38AvTO7LZPvl/
JWToIC7ZKZrJ3gUwpWGF/zJQAJgudA2E4c1gpPCe71Co+etSJxmHH+HLQT7JOScG7srHClEPChAA
Nf9k4Di2Zzo3MfdVAhMTdov23HwnUljVi239HH7nnLgoQ3AOa0nvwLEgBsMA3iRyS2ZgP0/7ko7P
+GfSCUtijCshHKCZWzbM1bZ7DC/w9env26P1ZHzzZL8P/T/PzxC80cL21FAfSdN2hkkUAtUiW36S
R2zLPgcPFjzXmskxOE+LlvZBl3Za4bDZX+56vE6kCYoXuJ96ZLE/0CbW6gy2K4Nvrl7VyfXxsor5
nIgDxwdRdxBbQhaZg7lastFV8AVCsX7gcUY+UwnAERdQepjmAFFvkft/8HAINQpXej0DP735wHzI
xj8q/6j0t9uf6VpqGy8b2tjUUzRzZzoeMYRu/+LZ87AOl0ZzPbg0HGuKVm8wcZi4+56VLJ6GE1VT
LvD7BvE9Ipa4YLD7O03GuCPptiq5YYHMf6v5w3vt17gFKaCMcH0xbQJ4Nos0ACYqmCl6THu6WuHV
ICqq1ClBvLZDFm2iZdogXidpQm8KWE9an7MJ1FjKENeyzm9oQTZjjrgf39ny9TXHcYzlyH/w0Fdt
BCD0dxExgGqZROryvjmznNPhji7AsuquKgSPwWlO7AeVJI9V0fGiJ/0q73ZWFUi5pHbYY3mKafX/
XsZIESg4R5voHmEx39pcdclnVFBTdlxACW7TaSr11hq3MZ7q7AnPHYdimWwDDlKYAtcQBsIIvcUv
lUJqaeaB1MrNm8F+BGUsRyq8E4RSbK9v53oNEh5Xmxzg2BlKDmZHcIVvCdW9OBMruu8pLSJw1c8e
qHQpTJfDcJlpnEzklUOsBpg9rH1TBUsShBCtQaXXsUnyR0Cga0t4skb4EPixprA4BntOUObFXqsL
SmdRgtHhCy9u2bYwKAYCtqrOHskcWIFbSXzqHxWhNblWsRhvs6Pq49q+aenWaIXf4IgR+utxsr1l
q+B2U31WwTbaFzvhmlivIz7xGxfRN7gr+22+MzX1HX0Khq7PLdtP2JweQHGpJn8JbixkvAZYdgpJ
3cmb2SmdaMsD08iCZ9wKtlrOBs7aeC9bMGX1W5PwPpEdIJKs/pFJhbKZSws6nybr8AT5ky9RxFo0
UyM/YbF1aC4HWKTKfcgUu1wCOwneRmCWUqx6E5EZErPtB032i9qHZ/BjYCXZktB4mnQ+BVV+OULj
ZrGAcOgg2NCiS21yV03cYxp9znOwPsZQI3PNLbnos/Wi42UNNC52y8hr+iM2/DhsOS5vbZNdmqXI
5cwFeW1SnZ1rHC/N2BS7ZUFYgJHJwrMkr1pM18r9TI1XzF9h1tg23NhgnaAPWIy4XDoLoBQl6Who
/NfFQfpL3m+p2rLDsYcvozKpZMQMTceKkElAx9XTR1DqVjALYpZ+PqM7i/2fqzmJM/Qs49HQtuL4
CEtN6t11dKUlWiaPOrhgXcUJKyrGFWmVKvfQB7+7W+kcwQJ5JC37Jgp/H4NaFEWk8iB5LNzVx2h1
4Z4LyzO5pJN0JUfQUADmgCRwDKTCL+HoqLJBejn+rO3iwj6q4m7qUUAzMzF79JOJykZCulB1QjCe
NWZ5lY0LJetdDp84xBhwBpxYkmQAgsy1kQXAU4rT0+Ym9hEvr8AgEzWmXP8PBctpw1eYak9OZ9LS
Qoql+fzInnPpA51ojZ/daB4pZqW8C9wrmLTsTrKsWg4LciyNPoqlNEk4ZuNwKA0QHjqDXiK30RzP
MEGttEtVce9eT4xTmw1h+igHvBBJAevTB2ZwDJGKfoyc/Yuh353y1BHMduoS6+5CdMk7vH5p/UNR
vOSEIfHG/v9FFbrJ4AiSug1RqCgQoa2iT1re4rfmlj6Xg/as7Asx8cDK3cDqJ2kV/UebfUwLPxo+
T8uKNbR01vzM5YpdCxr2JLYXsNTFnSZasHTQv/Z1yPs+PeLEmJ9V/2SN8fljkyZCJIXvt/9v67MO
7Tsb+7SZTYFO8a4hJk5ufuxJDTu/O21StlkqPUvIeh/DfZduDadziFJCL+iFX9WsYeS9zjw1nKGK
wb5oS7m0uUofc5qeJbZQ9CP4U7XVIamJlj1jl+e2DtWY5K0MadBeSTE2JVS7cdQZDeHVjekyA+HW
SIXRZCba2ii+7cUK2dctpmEPgUVCDVHBitDHMWDS/qhFaHCTPqUzFCq6O7UC6N+e6/BK4+g1x0EH
RkycPhRyGOsfBaxbv6pK2VtGi6vaCoMrxoC+BuI/RpnTmnbH2+eJ7UL8SKYN/Btr9LnPaMxj/lRl
AzFKPcG4aNZ0QjkpmvIoZTK1YCc+tc0XRjrBu8TF0b2PlKC04c8fMeuE5etKxpiUDlHP3q4OLs1E
SThc/D2JM+h6dDebn3rOJdcI0AJ7aCsiyBWVtClE8DrMgyeaPc4sIWKVOXTS7SXPp447sYBByzyF
u/5ay+q5MlC4m2U2qSjljaeniF9Q8YxFK57BOWJvyadbqE2FhALuO00yWvlDJd/410ceXVr2bRyH
I4w3ytGO2gFYZOMJVcDI6iMPXqcl1t1wDYsz1x6Lnk4HlhFIdeDBA/wlzkGzxmlvGiN5K21rjYRz
++q2iuefDAcqaRaR5vAYmQKHtjNxYfvYggnjSFMTofvA32nFw+/TMj5kHJynPAI/wmlih7pyl9KA
clswijKxHLayICfOub+sse1vkbbsmSGRIPrdMGvDmyFxOmYkzn9YTPiSyhMp+zcMPB2adCDoXe33
Qv0pna6l4jq7sJ2GvjkpScFDc4QLTA4IQ1QbvY8CLA1YIwDDiKaXZchjfmx0fdm2cx43WkgNSFD+
kY7j7L4JOEcF8ETqrZdH7l668s8popQS7CHIe77BCaaTG43bdJ6RpiuJbCYFlWGvgvqMBcmwtiIb
JZmtQUFnLeZiUR/IiA7lpi3iVKOayZpOvRRt80w4J3S8ITAilZYvYRxSxq/26RGvMblJZ9iNrZNG
UqPOzNWHyv6pdgCjPrXwouEt2PS3AS0JyRy46V8BiT7LagXothxu/7ZbCrpGAdFucJhobnfVOvL2
40u6N/R4+W9/kBut/63aj/Z8IZdcpRQT4rWO7PGT4LQUzr5nY1/76uzo2Bxu0D7V46inp389J0Pr
vuMb8SJ1HVE9VqshJn7INwoX/Zuw6pTGjEJMxilQNuVMtzE/FDGl2H+aMmZxwg6HXaQuHo0hBnQ2
UpyJUSwsmGBFMq3DR0+j0JcHfUPd7dYYZYmxUGTKoXJ1GtgzPj+xuysPdsW3/oCvsXemBkA1E06K
QEXsXe/x6nazL26CiIYs6JjlgEM0UqPBLgg+H7Nl6rsISmRZ9FT/1jonzH3VThT/IPhVB8UI0Nv4
YS/NDAa1nk2W3Aqdwb4KEnSRY5sYOVkFQrVZYx6DgIAprSPJllhMUDDiB3rV7PCLFPYPaE65mUqj
3LYlzR2SCffPKImCoQRZHSH4UHkMmapJz0TnLZRA5CIbjZlNSI8OMRAoAgcXExEi1oiWtiWgBfzk
myPIQaSQskeG16q4K+7Sz1ibOrFSVrxSvzaec4rEIUHh2AnuEuSvVlr5d+BdFwqeCOvZtnbs5a5S
KRNotYy7bHAbMPzDyfvBzYbiN+1XGkLgKjufhOxA4pNGMdZ+PuONi4Sc+qUV+vvLyK96B+qe/d+x
Evgeaw6Zh+h9ME+1MyQVqFBUP4FpdzMJnnGGXerHLudcHQD4yDXBFC7znjAyqdh97zrKYWOkNJGT
zvqL68ZmvT9khDffDD2+nqUYTOA7uNZC+TFul1rN2uoLhFJhFojPDB4RVArfunO+BCaH9YnX5bzv
1ONxN+5vwLGjEoO9ngKS0I6pNXO4cGv9opilhn7BE054HCnBnihBQhSfHWwibv0iFekp2Py4ZLWc
RXkKD0GVMO3KpCxQK+ky9HFHDnS4PWHr0S/z+mZsz8obvsWl4WJegJU4oAWU2U2TXn+StLg7SMjg
UQ3yStFcjHY19p+2iofXb51JnkSsxS1Eo57gqWgML8DEyYIKDARSgb+St1vlnrlZhQXaInqjgrjZ
wsMhURZ8MA0ufWNvzTsL8uFRMlo5YcCW01ORvaCIRzu9WgmXcLhsyhWXGQEnecgqUofc1eA1Terh
DMntuAWW32f5oPRaCh3NbD2Njcps0BId1pW5aM1Y/wbRKF/derHghoA+iHqkvrXrgl6QTZ+S4r1m
i76BPxPsilLGr2pWV04pxtRu0DwhhAgPL6IH6mHybRxugf+tyF3eGf+TjIG7o8UFJJdYIejwXvK4
GOgcnSqxxwnHhrzHtPSXuTCYGL2qjL9qWY1S22SZSfYWTwX2V1oYNvTlw38/wYkVw7DQ/mM+f3dz
Np9O2J2TukTK9CXEe4ZC7x948ApS4rCp8xQ1NLWa0D1yK7Q6djbWB3iDU62YSju2EBQAyudCAF1K
FXqrtQMWASlRzvhls+ngMU3kDdq0YH5PTCUulSEyIrsGaVhPxCnOg+jts1nZJ25Wo1F2Bns9qMSJ
1ON2mMD0otdDlwnkRfTNv+BJETEjiEGY2zBMr2SlV1i6hI6CI1tAHKEbwXsFnoizNUYjMQEeY3UB
qGhJWFJP5DGDWwqxf5VY6mov5nrfx9dUx6jsHsi6ydADJrizDjNtGGWjP+590hMalTK5adXpCBNT
MsNrySEEEE3D3F4aUbNRz8rA58Yn1I3DDI3Ghy/VndnCpjkZifxY/ohBsm+2yJ5eC96O5XLq8pNU
t6I+5DGQc4UEBKWvoJK51cvvGP31S2P2s3PkZ7dD9TgffCv+BrK5qcf3lVtO/jhu+IgA84+Zsx7w
hBE6PlAQGRTEkwHf3I44MNJ9dtpI3d7sjPNP+s1uovTXBJTxqg7PkY7ww/8uTXHVVfL4NyUJ2mh1
HGfg4CtdZFFK5KHn8iHGPUBclVEU2Iojzvc42eZaKJQoly6C015qSCK1DSp2dWs9sKjDk6+HMlxG
R990mexexGH+1FvUtMYEZsBZgQTX5VHYpUItdny2hu0qS03LqgZTC2Pm6SHoKjKguNXDVL6wfAaY
yIwfenijweURHIX1CcQSG2DdIk4O1fnxJho8HrWzoU72GhqsEQRj48BYxQQ1q6h2hJCgBd+KAqk0
8/1ND41U0hx+kzCm+7FVCDIIm4A7x2MCIgpXXSTmndaCGC3LiHnNbpNOnmENxl8Rac8zYQ279USR
NEcR92R9StEu8LmpkawErIgRf50A3ubSj5gJcyZ4x0L1ZH3nmp9mZpq4bI9vhN+MlBA00++cj7h3
0lqSy2xyAJzpi8ClRYsW7tABXspRGOl4gxwfNNnG2njFqhIPbQGtIsomvqdwMUty3L/LK5gtIKWe
LosR+v1GcVp2r2j/mpIDac6H7XQ5aLnRkO3HAzXicN2U+CbWByj/TgZVPo6437LgCC6WOIqJFjTB
J19Yj/NVSfXlON9U/TPrgBuVoR0IJ9d2380jmeOOchTqj8fTVlxScYAYHPxJs+rBtTmrOiRZmMLd
b8skSNkgOvMobMlWtjvnzs+yL+jgOZ3Z8Sn1k0VQhFnmqAPVc8UGt2WqURzdEaXUbK+rd/glYob/
nNsdBf+kzCjYW63RkkWn3SqkQ5yi+xOCJacg4ZJIBsKvsNid9WQfNLsUGVSJFXrpu5cEOxblMEGM
yxgh/SMYaqdNbPnxW68gAl4hk6UY/e0zD/NJC42jpglqzEXBB6NCkzgyHABYm0EOxwsJV9/BJqPZ
yEPvY1arv4aR8saw70+VGEXg/DO/xVKvO8cu3wEdetjqUNBGDKZxFbdoj/i90ncFwYr0SYveHBtN
44PkCAvGj5XJzYpPzsMWFEidsc2ATGdMXSkw273GvmzYhGi7WSjM0d3/SF7ydAT9wBDajmNqbrB8
HbKIne3FTuP5V4BOuyM0UZNyI9niKfJgSKjE1LsM/4gd2xTuwGMbXhjGaXsZW9pk4Yb83yi9ReXC
g64nV6EL1vcOuXGoRd1em0HMfrO7k2SK+3cum6B9yTmzjClgkmGPwdIYshZmg54F7PVDjvCvkRIG
82TtupGXlxJe5u+V9varSB81N0+GbKrvv7sopLnF4KABjFla9ewrPacJcFTxRmDGVbhfanJ6keJk
HadmaHlEIgHRmpyGQ0qJhORorgfspyBXS0poCb1neUQKHDPEgwRiNUYSS1kRBpkS7uqNWsEqol2G
dVA7mPurXBevuWDLblZW+xzewf9cd0Kh9KhX2g5mqze+CmKuPppuClTdi07R4KqHn/H5vtXbemi5
JS8Q/yRcqLVKd0ZHmG71jQ447ECl5CS4r+TSOn3flY3sMzlcIrdKbDJBlErj7KAf/kjwguXvW/Bc
yEvYYbutPcT27Yrfl5VWixn0yriJ5EKG1fY7m6e4UEk5/OVl4vV+iGTWE8lfpVA+/b9QxDJaHpCC
Ot6pCqYT1zuwiP+lGDfwpmVLPDhIVsm+iCirnWtTwmbN4M7BuJFg7H7offIW/IFQ/yZ+iP36Tefv
O7MOtzr//zwNV21Uo52eQNxjm94w1f3MYjwJCnOWHkBYpPFe/iXZmBkmLF8TTtwBsPeiWKvJQR3B
bXAG4S8GeN/nX28+Uhc2l+7I+EfbRp/7RfFVyRepXE4lBUzzDAL3aus3Pky7NaVfY/JY8qzIcWMe
WmXNOUe0LFQEwNXQ4wJytCrG288KGkDXcj3w8XPKvmd1eQxp7F3IqpuUOMogTq1vDXt44rwb0s5E
bIoS32dwZAiyKlGQUqmB0gi/Gnr7gtJFjF5rug894yBsVFiR4r54jRNDyCn3P0sa9urXXi4GT06+
kj1mHDYjkKUP7i7EIg/oMBC6nfingZgrESevEUegjLhC9k6rAnXx/6CbKrK8kS2FSKuXeBMNkXHH
tp9csCnrIR9T0LwvovOx5+hJVnjisfpZnj5nI7Ftcg9ZJCyFUhpIVK086+7oG/rBA0/Ti+9aJUYK
G/i8MVD24hmvvBFsKbiDSY79jQZe9isyxNybkzqE4ROO3xVUCVu+bAwQL9CwAtjy2z027DU/Uofd
9tfCqVeIVm6+A49Mc93mBlw580GE13FVtX7K2pod+TUUhMIbwnDAyG8DPO9kE/hVtrqquC1k7zd4
Zu1edm+YyxMoPmA302pVPH7q6YbWwycD4uwED5myA9Q8lkyiNm83N/R3T/lbxSP7i/eQUAVzsTl6
wkXchBdlfyJeIBn3ZI1HBNZZ4/g12rU983a4xf5w3NhSwR/L4LooGnGgq9QEbWxy+SU+OZ3YT4WN
NT0ygLdo9cc6ffu67dPQX9RFsbnv/pgmKsRR9IPCIG+MSdbXfK4PdpWGFg01+Uiara3bs1G4OSKR
yhB+H6qGwAKwB/+xqFXwD64hVkLSvCKGW3vy7eeFzrHoyEtMxcejEcYrxwre8qJASOgwnzUMv+/O
mfdXJ+4sypuqm+H5tLquy7BZKaxOpCZVZ67wqbyY0utmF2HgAWzWp/H/j/HZj8NaXT5ueqOLL3H4
QHyF++/6trPN2GxmC2FpMye/CL4knHEeiVaiOJ2hTj40PdapNHKC2RhohKamwV82igFYYuleufjC
IOcIlFkHk0hEl/ZiVS/Wea0Qxvrz1eq4sMhFa8AbB3F2qKBllwr8uRxa7mSMdwtJ1YfNfYeSZbT5
jcBkyOKKjwBByV+9Ll4Jx/PjpWkHqkyWuVGy14XWbvtzvMxZUNMuKkNSr8Xg1TGo3bVZTsw4xYXG
cAsWst6wlxFoWkbGbkWIUv1Ytrdneq1Y8PlkEfqdua+y4Pszku8OuH8Xk/h1iA84l7f0Oe6hXFFk
Ii4xJJLEv39D2/J8m5EvRPsVoIRO93ZblPqT+8ojVurPQqC+mHJ0kulmOB/MlAkaHPOJ9R2U6SeF
0F7BD+TmGI5nq0Nox9Djw/Uef+mPyHsJSpVp9PtWRmFQrd983CL1EmEu+Qt79v0bSokwBtBBON9p
xTIZBaj3UE9/wuUxCmNeaODO5Vv6BTIPY6syD7OMivG6PC1PEBwrkAo9eutLcM4jbCQBUxr9lExt
RTqy2MYxgctktvN+cFfj2xyeJ7nwMuBjGQx0vw9rjx//MliyveJM0QuKj+MxGwkTdqBcDv5NdmoT
kimn33VKqY5vzWkq5LRFkHY2gIJ+tnT8FwJf9L9RsZo9aukqWHU5HVmqXKge6p1lEsMalUppzcT1
277RoyIkiJ9IXUIW0PuHFqRK7TYM9s/Uwz9xVUveeuEvN+/dAaFmBPAm7dMVseHHmAke/ujXTSBo
X1dsSZ5P34+bQj+VsgvSUcTD6TZOXmGLLybbRJe1nppZNH9/YXTWnuGe5Z/9xre8R062zqnDCaBO
uhreHKeZ5imjYBI6ZqG+iIlPWBPBxMjZ20YCi4vL5PkVfdkgnc34WndxA6VFuSO5D4sHEGpYYyD5
3dUVTVB2ujhvp1Fj3+yuun2Z0dntm0vsGZMwdJDwemjlMLdU+FZow/5qQVc36DuiLQO6l6Cv+m6u
/zTHKIjacY6AsYS1ku9D0X62ww9ZyCsb65ZzHNbiadGM6eYDcBFEi+5jssnOueUZKNLCGQNd8TON
9M0eAD2Z1l5MS/odZ+I2orbV86EiZeWzsui9Pz6mZ5w7T9B5+lJ+uCVnin2wdRvPXrVAQmkaOmBe
jTc+VRVKrer6nLa7NEJjwB98wkWA7/39udMG1CEQoKVRZ1JoCDMzeGNkhygp8oVuk4cCsK8dPQey
FrLU1zXGxuGojHYc8JD8JtKN/HdsuTIVFEAjyj3jA6fzti1W6NdFJIknuFmliPojkae/gVKTMFgN
SRzyyiu+XsjbCdq3rtuCw9BZ1xTMhO/0Y6AEiOExGD9Z1abRfNhmeSDlfZGoT4yqKgNKwzXGPRgY
2Pf+AeGqLmvMblPOmZ1WlLCVyF5uuW4L6pplYduV1v+HLLbtDOthV1z6COUMt/F9D2cyDTpyK2AM
82sp+NlmtipJ9ElPRmdYr1H2xZLFyeZZSa9rBAzUcZBRL0Qh9L4FgGCGewBTEVOEsu0cSltGPkTJ
f7lFEGC/3OHWFMuLRA3cZci2oBVYdEJ9q2OiJYPPJ0YqPaRDgn7LqEZGKlI1kYDKUXdnlUOBQtyh
PFVcP4Z32DO+rgZ67IlVSTxldNycl3KhQU5NqwAy+Nz0pVVx5DV2/ArnnbXdOrYnY/n5RmN3sfjZ
dfzzM5nMWDBQRRaAQ8/7bYMP/ZivC05qKWeAiJJh4Qp78vfcgHkZt05UtHX3xRlRDjohVBK0UNhY
M7efHNvjswd4LB5QnAuhGUx60VgLo8cCR4/scpGY0P9TKX3zW/hqO4XV6nLeZgKBK/GmsvJ0HGZZ
YvbXBFhRe1TZKL4NrlkBrwCPau9d1HVD+IBIlEwKXhIUorTda45iGnO3PdyVi1P7P6E5oafeO5vR
KMw7N0DwGITwMN7dbDl2yhn3eNPQz4xIQlQNq8OYlTaz0ZnKIdv2eYolYQsnl8h7Dn9N7rMfF73r
7glDY0yCl6RzWRga8dHqMLmAWjTL87khlry3DfdgVBtwwqohtebfD/rdbPZDJ+vteg2/B/WJAeJa
Gw0c7kOs2Dpa5nIT1cG/arYXkMSl2j9xmMvKAvkv3KKM0giuJHuzB+Bl18cgQbSj8Fxuy+xHBkhm
RezbqU1czDfOQzBwvQ5Wa3B/fj7S3QdmtB1Ad1XMCbaLZm5cEfVlfK27ew3x0Wix5Q4d66ku2m05
NzyaILa5wdcjTOBo3vl3mbH49wGenPypNStLNDe0fhBN2/u6rOqVZR+DSg8H+J0Gs7rEXv1o+bVC
3iF/y4OrLYHYWhy6pg7yaHbEoq2+EEa1WWon31uYHp3qe3C2MTGM+V47fu5xOwU2ciuuR1DobSXS
nm2Hl4bL9mkmlf+xhYXrZL1B7AfnlS78YdsGbCOpyEX4CEykXXfs4GLDHvC6atm/EiItfeoArstv
ynFjW5ouua4bH78edB97POuuQkyFcqDvChotngPaL8bvCzwRuPUt/7aOhklv8y2QwRpijTsoUSgU
N3QTnCCR3YdKO/v94Ui4LvzolK9cXewEY09Ts/7FDS8o85bc7SFTvgV3zqlLSfU2W0cxs/LaZyek
EO5Zd57JsYHpX4VGaqAqdGda5uamtrl8TfuJRQIPbcA+9/7Eq3CJYRTf2Y0t/fB4BZ8ip6tI86Qb
GTBsFnBOBhC43cgdtMRiDeCXfeMAVys2r7498qnsIztFB3dxhf6ICVbyQPY9qtthsyoN6nebtED9
0iHwsm7x1Nk+sBLBMrl2DMeZMKx7ipqUrEnndnwALyEmJROGFCNe9J+Jufhxbnp4Nv6TzpaFgZOi
R1wMP/TkkaIOTRU5LTKLIR9s7wO/mW2ng1asXuSc4QQu6ofTcSvt5BStbuoMcIBcPDjzAbPKg860
/0rRv8yPtpxiJ490TkcH99gwUAkpi8SIH8C2b+d8yhaOF6mRRmMQriU+zpfl4zyfYG8e6JwnzB+F
AF4snYenGqpPcznD0wYIXa+FnzSZFR3v9L6EbwWNNAnFQ/fZRQvA26cZObrS67JyV/Ots8ii7Ki8
aysQir0EwWGm/UxzYWIsIj0TazWKwR31q6BCjeWOeerayckb3nrVb+4ui0k7gnxnm3a0M54UlCpP
+cuJ9+MMLKx0hMBITvcfYD0wgpbEPtF6nRjH+436+m0DTF3L7Qhp7Kt5N7/1U1GkbO/lpjlHMbZp
+JsvWE5+NnkTnYSIG+8MNN12Pyc6usyoVHwBDSwj3EkChXq2ac+6sqAGPjyJQUErPJVpBOGnbtTG
TeoaQX3mJT3u/qgYri74gThaRbJe3awbnFVbVSxlB1+nzjbGiLyEkO3vRmgBtw/nPpt5wYjPzftT
pR9AGKaxll+w89j8StIkdHeOXJ9mFUM0os+t8n79U63nGUDo9KO1YcrW/VEkbLTJh/Vj+J7fNK9Z
v9SLggRu2PZfo6Bge375PUtzdqDmUQ75kANSUt+IHDiyTij3XqGsEjpP3QjdJDL22Yx6YCQy0we6
Xeyw4mAL0wnCrXy/JV353e4WEuQNxlYVrvK3PU5z7aFfyzbYqR74H1eg194/mSpEO4+W+lrFU3Y6
zf71OseXSKzq2d7nqklcvyXOja0wHZp0U9uyw9Cg3ZhPLu7j15aEAqKuCFV55U+nuNa9iUWew3l7
gal83JUg322Slbgj133656aBRkRRLwYWV/V14bWSiesCO2/hYojQQgwfVQzLUXFPL1zStCRG5k8c
x7SrgVlXnrqNujif/cs4dSpS9juSTTr7PIRxuMazGgXlysRE1omVvOaNfTuiPYiHcNdD+ZMgt+lq
4N8mk98rSIhLHZIG6fTDLgdlM9ou1UfFsGIil70PJjhrXqDM1wEeYijXQkYPLtP1R8aMptSVMPLp
jOPzt7ZZa1mI6xtUzS0AGlg209YN+RR6YdKoIPbK6Nq84GuyoaBB1v7HRJeIQYuC/yYrtYYoSAVh
6x7pZ/jX8oxKlOmg8SFFC2qMDXwMBYDrAImPtOZwaGG/wgAasooQ4lpdwumO3JYvqaVgBjFSDE2E
X+W4Wvo70qy1IUQRJA7JA9eOXiFH/glTy4Ma148AvzO60ShCyHuLrrsMTzrMR4f/H0CICc3/kAJ2
DeBwPJfKnMggBNCduTdNpofar8mNTK0Dn60MDk5HOEiY44lMhl/EkGCbjJRcay1tQLXb+xdM+Nqe
wOPa/mivA3ni3iVtQrbkziaIm0ns382Bbc7tJ9a2rGwIE/bm2xByHgU6OlUyx1gYcqb5X81LrISN
BM+8NiYDqNxgD+XtXbBz3JkN4QCH2b8jrV/Ao5z8fv70G+b5qSz8z3yWe0SdlEp0jLHsoClCcLni
V1RJ54cYKrMyjDTJ6/DD1q/TGTInlB8bK/2yAey9J9fkyRXs62OaLOnfiVHgbWeg4zPF0cSPnKDV
6xdROtHWNty/YT0O6Yycn/a/A6MfaF89CPScnD5nhprBUyw1TzbWSAqlIbAuybt9WFNDywifB/YI
4mmdteoNokTvdHBfOSkeI6aOUSgsjFfdcHXeR0SlKTuOlQ/WG3Ypbxoo8qnhhGtge50kcT+UVBj3
ltc1L+2X2rbrTeBHj3dqC47/mM2ObceLpB0PrYFgOV3rOgOr0pXoAjJE7VM6sZML8tfMowVZENe1
A+J6bmW9bQX5+BZAYi0JPWKnPN5tqy1a91qTAQVOZCV5gM18SY16oGRtOFTofYmhtIE1GPTrBvKa
M+9oEgj9+Rcu9U+1DPWeZKe83DUp8opub/C3Lqune2Fw5sYMhtKmLMkfFPceaDhpld3eF24PpIYt
7ifGMxU03pM/tQFF6I1997MtWaiJu4zfgPLK7OIEhBeJJLOIAO4Jox7Tw7CScmkOfvwdKr2Jzv5f
SLdAnG3zqoKAEvViNRx5VYV55sEqQGeNNeC25ABi04njB2s2Z6CArqlS3ENDrfbUDtM4zrhH/+VK
60yE4oZk7zq350E0L0eLu9VTaNjg+I7OsIRJXeVqkAGVIrRc26Ji3oevvI3xGVeeOEvZbST7EdYf
my+M8ssONF5XJAaRi3JGrFYXJ1qNU/YO8TuX4F3cHgIdGeCWvpwrWYfdFpXa/2npU/z8mTiIBZUj
JWwFIx66QhYG3mcx2Da0UylKKUi5jGpLs5zJNVGr5PKlEyfnm8Hq6QwaifUpJUmfafoAQ2QBXXYl
aOPlnArt86ro+MFIgUnZZRLYE0tIiHe0iND85cVKKo0Q5orPwS7m99R176AoGFKfL8gPAsI1O1YW
gafoiHByMLTZt0fLcgCAplexDiV5Ryi5JvUyDo2VuKXv4F0iXg56PEyF2yDI7qtER4zZcyQ1/f70
vUvu9iZSiBpMZHS02/v1LIjXgenJpQeTzjn55hhKaEpytAYLQJXPZViFzNATdbpISj2fsqUhtlrO
Yy5qVli6B3lJZ08D/mvRFF5dtktkDYCXPpedkD8PSlpXNcpO0lb5ER/UD1VrWe7TV0OJVrOlBZ7o
AqrStkRwUzazWSUKvksqQD9uUDAROC9ObFbxvCDyi6t+DHpwBiwOdo+Ycg26VXtLV4YTYIEghpCM
DGoi+EqZT2rYRjAD9Ausy4j1cU9jEt7BRBBHuiywOQdyyT9agZd3JzcSeKHDtnRtNhzdS+OHdunz
PyYU42u7DM8m6xqUTSzUi2i60G8NYBc5DeH4BTSSbxc68KXyhxlF83zbCcfd6K0c+y8p6YyL6EDG
yCq8mQ5UOYBv5DNb6SxE2EOe6QRGbMdgDLXXmf1AKorSasQg2BFEK63r58+6UGWnp94amcK3nNHx
WEhjI6Ij02dvS/qNp9XQILkehquebXXN7vBf1Wrc5TIupZRua8hm4Hx0YuF/e32mCVgM7sEp0wFO
RxNiOl3G0/cCpOI9GBKqDaXU/KJQ6eNuKyEL0QPS7cW2h4hk+vgGudORiOh7TBeeo9RBSWDsm2Jo
PVWhCixEh7J2EvwDH8wAZ4Qzb5G+FZYRda4xsG3lpy6XGGDWXhXHt0dWAQpM4shQqtxp7qNZFKMS
9XGDui3MjEQVGLQIcdboEOqAoAT0I4pR/sHd/jG3iUcdu7dUq9AZosUFONkX1hcvgN9Gawv0C6RC
q6//iq7BD/l9iQXE76ROz7uq3dPVAILu8njUn+Zr4XFhfd46qoxUVi1YcV2+yPf43y6o5NVINbP1
OXgIHlVyUPQgJtjAkx2QbdOBrjh2+T0MmJ6UkMJMj+C3UdzUfyMFyzdsiVrEdSdLtzhjfYejxbO6
Bxy0BZ8eaUCtsmf4qBOXmXsoriLUYKsBdAI372KJabR3WKMyRoDOYTq9kViELMCytN/zG1Q67NN2
5KlitEzPiNsGyrBx/OrqYapiqQ/CXkOW97Zsf8PS35jClkNo9vL9U+rhFz646ark0X7K/FkGyBH0
TwPcwXVvpWF8nXLfW6sSGIhpBXklnN3wA+ie1fTJVeujSRVwa1OdGF4t7D/S0Mj21sWMAmVMF8Xm
18+vrvMhrCap50bn66GD3PDAE9qcXAYXZX+rRgfTw6bZ00gPIEf6P9z52lWw+exTbRGolIJM3LRF
8XD+i9uQl12Eqn83KNJIr5e8LHAmEw+WQGCejXkze2tUfBOC+niZZ7vrCH1wVYxQi+uQnsQsKdNo
DVMWjHVMkMQIXXjmdlF/pS2SWeLjLg3Ek5b6GwIU3ZJsa2DWXX/oTe+1N01nL0G5XayPKFDS3a9N
rQ2pehq1RZkxfaJfYFQjN2PeyUbBj7KumyNkS5usKMN5CX8i6uAVkZ+ZQn2C+616n/RNoiTD7sFI
H4+HmwHxBOhE93EnZoFzZCdyUhzoKPpexrPlMBCDJkDD/bP22EK5JkFlT64NFCtedrUDxW3YUmpl
28NbW9hMo3h8FCJKaoZhSnFVwsKxg3/vJqjMO4dalqXwp7VvF6WKBBhFdFBTaOC3T69p8rFC6BdT
+orePD0zn/hHfbkqL+FApkrPgCgOuCpbOxyG3gcKT76f6t9FK6rzSv7ThpRxo3hrKVd/u1+GazyL
qLYeQ6cuhmE4BkWqbIWEIA8przOKNgPOY0fyWPU1FEEKjOYbUPDQKsKgZZHv1NllxmyRjfrOMlgl
9G4qtjZCTi/d8EFYoo/i9km0ZOuFKVXuEQKEM4HYN2m6/HwHIS6n69KE8v3FacQ7or/tVvB3XNrJ
CD40iaEcuVfzhHwPSqDX++FK8vx+31ihW6oTqncDd6UC+PbKxsqgrO/bUm4vCRuiEfoSZp1MlVs+
aso03cFu2SQJLZNHGkkkLxjksuL/pz86bh4LW9giaHz7WDsg6b0Ax8spI/sEvCDs79q5da4oI0Nu
Df3oF2HIItYmI/Ccn/iVnvcaBJfDVqBzDdVEy89TTVzS0g4wFEIWJSXoij8BsRZUDe4QRQw8xZ89
uoF2G0mchny+HTjDeqCmO0eQhK5Z7mEPM2JHeR4diVBBACOtmCBktwPh8zOESEfQNNJ8NfljvMSa
RS8SuVqSfHWhGIlIoSyQ0rgPsDgmx5ESJdakELewlBBgXCX0r4kfzy9dkBD5/w6T+PTR63EYrbMy
chBdzVgxA/S+FPCoFnJ0+XAVLWK1b7P+y9EES/BMe9uZsk+WWrKhZHWOOZGJNCIVYi6gpjNE/n1w
qbBFcfWgrrTfhTLElbxugQwoi7t9tfQ6eqCF1Iq4nrHBPUtmOdQUIu7yNapFniWBM4VVjRpmEwkK
NY0JP9YIgVgvv07bQiDD+7E551RQbQQoEwh8FWahHuX9y9aITgls61Jg4zARBVBrPCyK5v8/mVO/
2Rn76IgTFSt9PJ/APc2w6rbBBUrPJVrh+23AG2vOA1FR0EJXApg2o+xTazGhY8sSPF3vA1bd5TNj
/w3L5uOWJ+UB4rRqI7h6mj7DkKoMyX9sggBs4mAnagO54AJFuwg+KgN2E4W4IK0Ap9H8qppUCJUs
r7ZOgd5mYR6RcqNQTSPzKhh3V1o33pWpU8Hc9ok6AzUTL0cy1Vay61D0pnqrc9xOQJkU5yt+MD22
D/AmxiUc+H1pvKyP4AP+YxQRLH3gEH61zh0Zsu4Emq1JaQIq5AUnmQ+QJAl+KsXp9UyGV1dDOBVg
uWHBr7K1Lf3wh9Z0V1/eeZEEIsITQRHKaJH+Krzr1k/E7QT9ANs3T7zopjEnMIX/X+7g98yrjzD0
Q9zuDKqDPItmlAahspRT3KRouDvQNsMiFzlGQfLKSIxijVv7gf8WvMHnDvF0U6gZUQMuRSbtq3bL
uvd1RjR1+BnxIAyF3eZMNa7xXKawYqI0wawK6eVrTMrGlzfYPHHmvWTirDstiR7r4T3ACgxP6ZO3
jQjF5BJ8Q5aLN5+AIPbXjR7v7sn5TcFzLSeT69b9x5zGTOcdXQQxazgwEZUrqEEoziZhnb/P8jlD
Xw/LkOtyWKS788chlCQqMMsbxTmibvVjowAX1wFpIKfu7LxrRQHX4LM5gMWCaSgPC5fzdgtQWOKi
kiIKFKY/cDr0FOKmbGeWrcWGlo7ABesNHJxuDOiurdvxHawREM21sN8tloiFiKejOYpQsCSWIJq7
/V/bwNrY/pKqy49gtJnLUQAxikLHvaCdsQgLSUrmeggyrtRCzNDfC3beZlgXYL3W52f6pX+0SOqe
hzEg3JVo8MV1LX4fm/TeDPF0B+ZagCo/z8yfmzT434MgBI/rzlcXui55o9x33Wg5NpKZqUYEZi2Z
w0cGPuAsUW4AVZvVuJW0JnugOJo/DOY+yppsBByW3DA5L7Q5vroazVwyq9gNRTEX5XRZIFGzoImC
bYeXQI6VlDN6Of8xvveKoQHGQ5gcyvHKc6ggnhzWaaMgxSCFtmxa3z+QBWS2CXA2u4YjTVC36lvb
l4Zyas6Bp59xRzydLsKY1RnRDRPx3Qujtjtp2yV7V8wYo6MQTYB0wJpbTocq2yNjllNYUJDgWBG1
AjedcstbEXPkWbvgdco5ClzFUUDXy3Hb8aSSHXxnTEMqgTDsjIbzlv1rRrGGQf7ySEYRqXagmhoK
d7xINaKANWZHkzj5fCIp25JQfPoxwx04InWr9AsbkH17ihuharGD5ckq5KH3bVqwxxoRKsYm8ZJE
SBv57uqSxmRJ6pH9/cKUxnKJ3dz5V3i/2ECaoyCZNZfwAx1eBZxf2++HDnA+LUzb79cxGNG2z9Y0
VH5H2/4YtEJIfo1ThkjvTgE7vA480bl0cv0of3kuzDNG7ifdOxxnDzg2Sq4UIhobKquZmonop/3j
uIZnrlgB02mbr+Di1qFny75Cai3iXn57yq7Kf4Wjxniue8osMuOKs7tCMmXuw9+8BS43L9LxVbGe
XMBijjxwQ61GDcHoF3mSz3m58QprDRSyJNVAKZLkA0oaa/NOmxRVhZTrs+KHDdVr/pbKJAjxyz1C
asIVabjP41A5A7yNZrTRrDidu57QdSgvULj6u+n7qMhnRrFo6E7DHaSUAp4241Tkk+03742iSVHz
BF1BS8cIH/eDc8zDzHcTcJiKv+qONCMl9kiH36EQ5fXbU9vGoY5zR/pBu/kx1AJz2dRozYTJ4Rl3
0ukJsuLIb+JBP1rtBb0IyNeuoPTJQByg7Oygopk+HFMiqmAmNDG55l+PydB0TNVOtVRglchN1qTH
Es3d416wePjuqS/jzErACgaYHbwcZTt2rKHg1d9syOQVFHHXka/J6sVTzMNW/xZkco6MInXQ7pnK
H/oRgcWmXhXdRftoUb7bwdh+pNsIXZf+tUlibNbPr+UAZYXUwQTbx+rT0IiGGxEzUQDfheoTHl4v
Fjw7Va9Qmx90yjFv0UjCC0ejTc4DrPkfiU7kjs76bWQVVhYNi4S6QvBsjTU8dJamDc2TYvwApwR2
OYNNAGaTETtU7FtJkinwipmX2H9Drz3PzmeYB/lDzQ2WFCwVMAvxSBb7pKyo4e4WK1Uq48Kb4kjE
zHAFCU0PPtaq9Eo6xml5/qsTsboVbmbETbKgU6j8jLR/G39Nk9izUxE9u59AuiTl4PLuFdeloj/J
ypQOl/oi5+xrTnNgbeAXOTeM/6BMDT+il5QY7/ljxoAlHJT8Qnc7tr7GqEIoxNV2wQgBevsIX1Vl
SdYByjJCon8DcgaGKtVmUCgKNKn7AHFy3RN+aBTj43yrpkmd2c/3KzU8Z0By/K+DsU113iud51Uo
gGIePDolQIAQzfh7WInWRQ92SMzP28phW+UtEOEe89lRdiEl0tV/t877Qz304/o09ejy75jIwsUD
MTH9EfOTfsD3KQOY8MY/55A3ZiK5V5M0LrGDiki2rri5USPuq/0ZGMJ933oPUY0HcMw2QOeXm/kX
BNd+kuulDS0C1h9DA3u4Hafgeph0QGXUEsVG56oSICXb+UgrUWLsL1dND/jx2PTHU5JYkpmr1hVy
uts8XSWBKy+Vxus+kp/L6/Ft9dvSe6luvnAJgQ97SsAkWSAnaN9+KRdK0H3Co73kVxxfnYB5Xd5P
Gg/yVnFT+43xM/o9E5TKEgpvN/QRDKThxQW/0LoGRuKQhgijJmQ6vEsMue06+x6dzAJAgLpCsHD2
kn6+VkpF26vTSnC//NV1cQlIfzFKd2Lj/bQR5D1keXghNB5bDnWg4lE8Smx7VluD2FWXnRDute2q
h4RzHFGfid4O5Xl8zxr2NyARFm44xTVdpgt6aEVMrvnpQR7XvqwERb2b/Fe3xz6tawG/YfLlyDPH
2fN2dtbSlNrmv6VdVEZI/X/kjAw0tA5GlwVd7Sv0XsW7daAkYOLGdJsciwOxBXWESxIAl1p1BnZu
2aaC7FvcQ4FRy7QMxykihd8K7jJFMDPUwBrx6ep/m53HG0tnvppqQVlgta5+6+BxebVKGOAUvIif
YtKQKEDeRtyUbZTIBkDjr01dv7pz7PpImoQjV7cAiqNJ9UaLPLPnMyaNtkI/oNjyWxtXWzrpDQH3
KFcA2MWlu6IcNpv4TiNSQQENT8Zlv6wpGYqCYruusl4hrzGpwIacq8RP0HifE7a0J0eBAcUhPW+l
QcEU1ImgyelMsIy/+Cn1jWZcXRfuF0B4W1wELquqWNgiuJkbspRJtS9ofrmUY4CJE56A8iYMd0p1
6yqV8+e6ufPLhTZHxEN5pEQFmwN/QQIEFrnEgEOTJ4eJ6eL0UYmTw0m3GyVCf0oH673mqRvSLnTK
MJHpMujF+g+OyOq59tLtJrr3RTsx9BsCtiqsFzC+T+gBk0eifdM0z9CyWuVUWhI+8VboYfmyRmTY
x2TriZg+XIeb0C7UFye7/9Tscyo8ey81IRdRq/kK90hy3tnMCjv32apXI6DLKppJkNRs8U9mjnhy
6QOP7H+DTSQE0JEgClPhuBRazieYpuf6o1vjLZRZcHf1EhaMRL+s8sJ/IyNbH0bKUdRWqxhquorJ
vMtzZaw4C4Xc6UEJoa872R5W/EcwJyOt8KiqfywTE+LugaieK9DaxpIavbJimCjknj9iuH7hv4oK
MOkiycdbir29dfsDF0gX4BMaeYtdx5vJ3xG7o8HD6XCiKkGIv4Dn7R10+ztD+RmB1QqtzdSDoKZL
/gEP/RBp4RnwpTgB8pZ+2GrWnhw4/lPFFzQE3Tg7XaLPtnspluODCZckfReCleoVKwY4v+NU1bRB
pLUypWRjrquyoo8yLFoN7PZiXzDrO4SyJsnLvMM605ct5tmBN707Kh5emjM/m7YRMZPfBqXhc9TA
sxCdXw5+YUHpf+i65thdGNID6rctYst04JSTz72jggYbY0JDIB/mJpGg10ybV54vPpTQj29jxjuI
zrW57p9hQ8Ll3udfPq83DlZiE6txJjPfg/eoL6lwSkemEqy/YrwWGreXWZadtRfqMrbrE0L4YUQu
fvmqGmQ6zO5FeQyBE8LSWzlGZjaeewLNU32NltoJAuYSoHfBpjOGpDkJnmBCdEqtF+iemUfeM/C8
WckQjuh6lUlr6jFi1TDYkVhDdRK5+VkPyVB7MSnY4blEQGxZ192uzAapjqzeSpPb8U+FVE11IRlK
gmDw0K/+Adlcw/phcOhIwkmI5jaUnrgcwnoISRAMWrdY2BUBBgwldIyNVwqj7VpbHQUQPNFDB1vn
mO7sjb/lxkyT5OkCH9ByCcyacFXkGrIP8rSMSGBQ94Baf5pussUDrxX6sF0SSOtCRuKI3TnWWzSF
/C7faTXX98EPwIJI5lU1M8QGzR9XvlJRXMWMDSHfxlzCyE09MVitFGlHuXWRloi2GQs4re46GRsY
lTK/a8HpvUnsYCfSNB+KAkEUbBEZDXgDqQhClEspOxTWNFFzZEDu63mr/p/5DOBGld9ItiiwDBZ0
rNn10POOOrI8WG2F7kdeP/FQYQuctuyzvpr4Cve/POAh4SgZuiHpR/hNvhu8khsCsU8IuGhmFw6C
a84YE6BEYMRl4fubCLtOCJCu0dilESGXGDSX0YKR/VeK0Blj8QCjBgGttCdJDWOD42Tk5Er7FYvW
vbwB7HYgw4XCYK0pwrj0dfbZgNk6G/zM0PBQdz4Jj+7AXT6/dPbHt0NUA/aZPDTLI+kA3XTi1Jeh
oB/EY+cbWVlHi69g3ltXV9yANc6B33OVy0OkokNGy2AP214b09BRzQYCRnHDji/fZSvNXV78TFSS
jsycbxbIuDF2waAGp8mGldfMQfNOZ/vRgPoBBQhAcAUkD2Gxvd+AtbcipsoD3P8lEyAzzz/XIjVg
/uG0s3dsCepYAsTHSp8aukFNjR3xkXnUYNj+pReI2pHgiXI390++hdFeFM7yRmjn6krzQ1hGmbCN
z3mtJp9prQeYh6NmsmldF+PIKXOhQXuVU8gbuxxnj83MYZpxMi0tlBGcSUQgnf8/vu5tgsUo4IHR
rso6qIetSvRDobC14pQdCSUiu/oU8rIaApIMKs7P9oDo5YV37++PbpEMqIqJt7UYJC4BSjAhS1KA
nPntJA3LtsX/q+X+bGlxo3Mc0ftuxw+P3YILDT4ibjLX+5vswsnbkdbWFHIKkovgXwG47VOaUz25
jOKFgWPma2CEHbHjHBfesepiJ6/A2Sj4el+u6M5Ob2jWdetXR1XGumqzd2JPrBcj7vbpfzJD+3T/
pBz/eWwHjvf6TlZ59JAg5KsPiIdu1tzRyp7w5Cqi4Oo0aJvFGMZnKxMxeUOd8JjfCskmPBzJP5de
Ibjvb5Owsr89vQdR9Bt4j4FA9wnZ2+GHQEoB4PNBYK2nAM0okJFSg0KephNQUW1seghR/FevHs0W
YszauAGQ3HqdGg1d9/WJpPUnbFiql90LBo5FIyvfB72kgoBTsxcxshY6rELQEer82UtWFWLaVuxQ
j6iFJcEKQOB0Q6j/4/FUYvRCcPSUvP37+uMepbxyFFgACcOiYf8EZOPRMcNNzM3bIfja+eyMCu3J
2J4j/9Us3wYbr0FHP/0dyVrigIFQvGKcCicXHkZm4Iq9L6nsJu+uqU19Q685z5AztocwRAwhkf1x
B1lMeCzL1/Nz0ZaUh0KAXsk73lf7kxOcGa9XOfJKb1yTeSMXablTHHMaT7b0slfDBlyg28JSyfAN
E2qQcdcynPRcx5g3AX2ePxsvVcrsfuhVd231FZQg4R6AihojNjD9605BfLJz9Fl0evba+xLIPUZC
nw9CZ1GLgV2ajAxMAwm3zRE+P9l8b2e0jq454tRkb8k353yzhVKCxM7Vbkn5iG+Cj7xPR6CwxG66
wdljuB3no3Xp6iw1HjPWgnju68J/TSeyzhqNDIM8BK68d6z2KY0lYOCHuI3c/uD/yiK+PHpPIDRt
uv4RBFQslA3CAgmmgVXqm0oFdT+aQb+dEvXbytRC8ybbPYUnvTw8FbSdo25eIqt16HJXyLSAbJ2C
fCCkXfNOm7zldD3O1ODPRDXm46Kk/h+DiaiB/a90KPBXmNHs+H6gOsd6pgyRidUoMQyKKnEGitCu
CWWHvtjpslJi4MwKa7urbPG2CRBaU8VKlmABne/J+LjVBt9XYe9SA1hY2R87I4t99M1fZQ+4Q77N
kutqvf/MA1pjKB01m0+3LFFOvOxmCLBwHRPIwTmhsSZ/NG1FfGiIFEuvm/wIUKe+5+5iRzmP5qJ1
zR7/qpzBI1lwtzZYs+GQ0r1ObgP1nc7a2ZUKfLisdefo/Bu+VSt4r7o15+gijXAVjbfU1Z7A7MZY
SyeCoMhZm+jWXk6CQ8JCk//AR9zS1kLS1zrsHZpZrGtQ/qgHinbdxrmvrQ7/uXqmJ+fdf/a0j/FJ
sp+Ei1kUdWYXvWn0RpI2udE+uA7ut4f82VhJfEXs9s94NQpYsXJE6Jr72lAsaAy56QpBGJOwzu3P
4cvwPayz9DLNLoAv3qcjB6BcQ/dwbht/2or4O2DQGKpVVgnbsk00lSdX2FSPMVrjfsMUanDNW7GI
jQ5fT6Bzxw0ob5VTWC5Xnc2vlKHo06ZRFZDRXKd77wj8KkxkF4PPMMiJOcwI0tQ48WqAAcptc8sc
lOQTA9Wss1/DDSPC1yaD6nkVAHRuE95Wq4TZaNEpvQIiBTv3jcO2XNklH+UYrQBpNZgH0M2Yh8h4
3LGBbz+aHnr350dU/u5WLPmDiNhuZ8tDrZSYa57U6J6xpnB7JZY6QxidnBwHSPsTlL/aog07OhN6
goyOcJ2eb+pTriHoRlXMP/TkHNV5sV61hkXzNYBzlhj9A7DytS1r7GYZdDfQQM4O3l3GkFIJMubZ
/V5s10ANeH7q3d0e32UMy56J5bJBgUG/ZmhO7mDxDyydr++/FQse0IqVcDRhYGfnbUtpZwho5col
IKC+RwHJAcZ1cNdwIeedjCohMJZ82LjZPQJmKuKuuz6O0yzorOgQOBPtXsMfy5A56koZXqWTeI5w
yzRcjphEEJTa+94gpLBbHUGe7z3l3OItoxd9HeZCTc0lFbtPRRj190+zh7gMmrui8XRpRDSVoOiL
/eA6jWbUGsPwtxu2SrZCOiG9RSJSJrQAU26XWMOetf7joTG4N9v9NjQlQkoh4kggtPR7xlkGm2IV
bKpdBvo3QYec5hZD0Chb2GQrNtsX0BFdlr22dISWNtT1PzpE/7NyOGOjbYT2xD/xFlIBDW8m0odS
d8AAelzEQ3/jpwt1ock/6Ryre3vUiKDDIzaJ38Z0nDhZA+QPoBCmG5c/88RziKyyHwe5P5vs8RkR
wukV1HIdZ/UL1gafgkKi+/GXXulGsUL1aBeTACpCAo4pkzZgibW3KDqLVtTbs6xabeakfXpdp3v3
YzL6l4sbLWLyVbAiHBdJ3C0sK7AznksGng0ZjGYhVROHuG7yYow9udX+NFkYNzCWDK3tUtd1TJIp
Vd3mt+SveQpoeHTOHJm0x8UUD5f6+avexbEwYbDxm7QDmgTFGx/qL4tqigc2/hGPi+heg1xSEB2w
zpfKAmjnLfVPWvVecFHPT7pB00vgTC/59EwSFEFFYPdzgRl7TfnhBmAzTEht+2v5WTnL/GvHe6TI
iGmW3RRzIGg+1f49KFAyludsKDdbO/dukQ5dawZ1xqIxuAnREWEayRYRJBhr9M8p9Xu9JViYVtu0
VgykoMcXHKHlC6y9gCkW1DLdum1wJMPa+kokOY43ZCQly4lq9aW7s+sOkh8Z5QhjgJG1R5Gv6N1N
Lokls1eVlM/WLTLIH3I4QzdrWTgzICBPKxZaDwtmUtiAwwZJYr5vP/o48EDSsfDb2QN2D/AhdikL
Rw9wbbvdYJTH7Z2kw2KT6ie52CCxTkFO0pI7QhQCKYDJfcCcNLbUCaRKJ1mp0V5qEh4owzR397OO
2yoxZBsSbCiNE/t/Fx5sNXgcMSNECso+ueHkqiE6GSxX3X3cfluYzd/gVwd6vwhakIoiZmsa0g27
iAilUZWs8fIiQNgS4wBpsZqltrY5U7fMuu2fzxeP0fM/HBYjQMxZUs4KF9o1zjUz8dXst+GDKzak
Za86Jfzimo/5qabXNm0sfgKCfYZZWBaEDMkxYwDWlQB125eSOZMHAB+C6EheMpZNNNA9b4jFEnL/
76LFC1U53uKfgVuzE/02ufp3thVI68/OerWwFO9nTBo34c1kV24BXiS8S7wrJiOa2Hn3w9h7aLSB
CBqodAY5GanUZ8J3gtgIgmG6O7Fv9FLMQ0/e8p65si9VOQSO6bzjOk3KLgPl0WBsGp2b4vIG0Ho/
Fizqxmq9xeAI5jcgy8UA9Cb0aXwDDrVLsTfO2h5c5giYIBD4CxP8qHMI2xXrdPLnGO71PWDkWaJh
gFRX5oqJLzWnC9dSrmJSoVHHhdJnycYfHwbH40F7+XAKTYIsd5i86NDnVwzpMlWehg59x16DeTP0
adyxVr3iMFZBHtpA9aI7RMG1we3vR8L2CDYEIq+AytbqF3yzdageq2E5OOELXbSYfQ8scwiJgcei
e780knjlMlCJVLwA6tZrc5rJ3AR+uUqC4ca20UEs+MM3AJMvBPIKn66+P8tqFqsbKaHIOvTHyohh
XdwoGRBXm9o34vrcYXBJp79ShtOV16TCt0v/Oqk9Nq43fy8NckYmzrCKsAJbmRpN8+mEcITWZ7Em
WEyp7mqyNgxymwHd1TjKejEwKXmiLQgGm5i9b9j09+vYJZ7TJnrSyTUJi1TcgjclOCvSnXtg9Unc
4srPJnMVq7pEPyNHvhJEcFMSuX9a/HP8yGkDiFI2h7QTm5AUAMu89K1AGkoGeNlHgj+FPwXUv0s5
GetgxE34HbfolbWexmQZfx1L05304XezJZ6WSSTizY2s3aax5RKLZPFMa13ENjwlIIazpJM1KyD5
Fh+VR7xaANNWD5G49nqq1byhniWsARiFB7NrMAdkO7EjMu2xGN9ACAO4iuh+1yZrDnSexOD9w3fo
+sZBIcI2KbtBuNidglG+SHF64dKveUJCA02Gll1sCYZpNYLFLEoo1bWIBInRJCReJux9+YmmBi+q
ElINOzQ3Py51q+E/lhR57j3kthHpYaPsgBm8SEPosPttNCpVrhCg0APNuEy+2W/aYRglq4H+j4Mr
b7pYXThQJcVHzN+n734UO65mwr7RO2GBC6kAfY5RqM908Vw2K7yPCGgU1xpVJdmrmjfTWrtcwMUP
t+gF9sdUp9qb/8r1nh9hc8DhfcSc+aWGsO/QjOgRZ6opaFST9Vn+GJCoVQKFiiIQzTdbDjjKxsHM
iuYLQCsl+IWe87Bfk/Ncph219eNvy91bwobe0qD8bM37Vl4umxdD1UzXQX3YhsJI1/uUZ3+cAlwp
o+y4+XPwwAf5BmQmwiu2ygBKQC8h9vs/xDfaiw2ab3YggSQ2mQEXqRVcwBaMRoX9CmWQx33GC8ko
klmdthyRxZIFA4jgQeC1eN2wosw+UznjoGhYiCdXA4emxGH7S/ksXamiOQvM9RcJzS5kjt7IfP8W
LmSpJ6VvmwZaDa0Wl+KNzGExIa2D6Agq8xO+jzOyeN52G97+QGpkFjT7sna9ZgfF0gDMVZtdQkPh
9sKpZjG2XfeOrB8AqdowmvTmfMr+zfBJVSwzMn0VuEs+UgTqDDjvKwfUCYTQ021/k3ctcohGox7S
C2rDBGQZFUl6XB2JettTx/nqq3trPsypks8HUjXqJ5rPsiQorc5IkShk3YAIeXpvy/yYbgXcxn0t
b6Vn9gMWq1RSEbYF5dsF9GWJCG5u+Il5Ji+UN3Tmak4dcjjt8DOSWIaJY1mUQ1VNRAB7SFuh4Gz6
G2zGtGTTGPDz5BY+LzpgZt4JjixOTLhqbeQUaTF+I/Eovzc5tTWAH2VS7YRjfsc4kANglfy8RcGx
v/mUMIAC2LiaHMxuKGsGsMfe5tkHy8nQAuO1863x9DjK9ONay3nx94Pa0MXkkin0iN4IQ7nqUl8U
sbEAr5C5EK5B9gu1yjebii8DAZP/0Ta/4snoGa0wDOjbjsFWUihgGyKVS2qYbqix3bEVGGJXuAn1
ZH5EqQE6sl4RLqFos+rbU46VQcCv/ifYFVNcULJ50ORoME3Mj7BbN/Il758LUp5e0xjw/aohWLY3
8IsZszH170izVV9G43DzAlGSWsUPKIckBRiIIbXBbByOw5I5txZxRdzt02oSkd6ccc1K71jx6Vus
Swa9Vu22BdSt//RirA/Cnq2+9ByRXA+JBBElVcOM/H7luhc7AcPfo5qhBlMeD2OjfM0z0isnX4ci
LYnoorO5EpWgRdZFDapwSjsWHKcJHg8tPpS+jNm8KwKANi/zasOopBI5svEDAH3OWTBEt6evGFDI
drka+7u22j4wlBQ5tG5qiKcn88YA/UAQDLZ6l9VjdFcgjdVSGXSICgdFiw8tJzBi3uKuERwdcBCm
U+J+FDE5egGoHMjMySO9I5aQjEz8VYdNmDydYDJKXT0hzCVgPlexISM824kaOriP86PsnOyavGyD
Us4QcfqjEU+X6nE7Oiz3/Ko1dZNhd06tKoyazcqgdRWX/bzFwXdQf4El55I8VG9N9tynR/6GnhfD
749N8om6qa0M/pl3BeQKIvVmy+5afR/LgUBXzQ1qzDqxcQa5CwM+W5f+vFQ8ICXjVBGJdOX7WcXF
MHPlJMLfFh85/vghX2mwbyhjkJwM/F1+Wd352zSwVPnWcRFRa9z2a5F+zSfw6UyBikus96fDY9wN
b0kXgSfJ9If5T5QOF4QFxsXCPO489DRnWGzClri/E3FUA5h+xhu+NK9qvmVaSQZmG1jLwYl6+Lbd
olNFa/iOIRfT6+f7Oe9aKwobG12JBGlBCxmjFjWQusP2HZ9GmGfm2OK1+2/1apgyVeMIljlcF8nY
mnl/iZ8sIErkpFcpqC3yv+3GTn1YgkMbI3HXwDpXlkvrukqqpuhvtFfXGbaeS2F5uGNtKIDRvB8T
YQS72btawqtsCRDlUwfEQw7qDuE/6+m9goAe8zmYyd6HNQ5yUGWwe6XQDG35PKwAEOsaOIQOgiLG
sPr27HffyFXqNJmbgL7CH4wiaAb1teQdUOtNkNRiV/ROFtUOzw3jDOusKSuMRNlFEOfxCOww+rv8
D5fHolqZiKCz8EmX57FXe4sJAtWEG2mX25W1QOFAPtNFZEeDegpyPkx8rmdXXYEHY25K+0Br0+VY
PKND9K/en/dTFqCAPUj2J16gb/CznjFBcXp5mM1MVkBT8axAXza/FAjZ+TICWNQ7pBjYb/on2EB8
bf+qQQGqVY79slpeSDareNuDYigDa5ZnQXofJw0y9ezYNqeUg34KbBRz9DNdrpa21WmmuE8+ubGa
w2Pt9rG42K6qAfLkgy70iXjvAR2gC1Cfpk5M/Jcv20yI/9uihtycgHP5660wDOggR4RdP58vBicS
ePdHgB4OZVi6B2Cu8EElqpfkTD9I4mqWPIXJ0hhsacM44Uu2qNEJcw0+zggSVex0BQuarmIyccZ5
UiOaM7ay0EGJDXMn4eXO3OkVx4mxACgbFf9gNwdLdGAJkhM6Dsz29ywUJDaRMuUXQQH5TUVZ8lym
PExWBpW9fMwJ3QrTOaaNSuWKmZrBfGBieFunB+lfPmKML+444AbdR4lRGNdEAr9dli7TOLImSnm0
6zXa1vIWuZXHChbYHepoj/qZ+0SFNHbNcy3r8z1fN86nbkxP8KmkHsxMYQDR3xOsiHuXNjmxgj7z
fDjd1FREt61hs1L2wGcjIpznzd2cPPZri8FKBY2AEQFlslUVwWZER2ZVtaibYL2eyH20FqJEi+Cx
9wHFstViYr6DBQ25YIwVEmx5dQ5OFu1SZNoRN5zrme4UjET+afdu0Lb8fi021FtkOT83TU/Pq6Kf
PfAMseS7J/vbglqjmh2Ym37jjbcq+aqDY15vdj8McYiEpOOr9Q3F5hWiYT5tpPrTVOGktE/mo92N
XHPt0W/Lx4fExgT7R20giiK8xRD3OoF6vnkHhJ1fsCgNPUpDNqZGVhLZYhQu43TxR86FghpF3ndC
lewKAvKDPJUqBW1nnuvXNsaZAc+nNnth7z6283egSFL8gee/Cugxlg606Eu9JUaqBDl7H4gFC+lc
hCxZJNIa2gOQwh54D0MCKPoSSGf9pkVjmFebZ1sWVFwDWj+tsj2X3ds2jg1/DvAN/mQduuIdPTbX
eD3jaw4X1ij46te7CDEymXYo7dtPCd2/p395UHJ4aX9qoP5VYZiXFD9Ir1ZHTAAId6Na9FvGvSNj
mYXPa1hLdC0mOnCQNXmGIS06kr+7rpHR7G2O2CJ1TdBxmjvKMJnj4HG6ZLS4J6ujM45CTuH010QE
SRQQ1STjqMrbIQGQY7FRLCL/zIBS3bKUT9j6t5ETmjCiF0Au/eeQHb0ZdYvCQit6nSFR+i6h0izX
l90EvI+U6/gHaL09ZIBsukNr0yu9Z9oauFift6KSJhqorbScKLdmSQe2dIcO4WyGK7GFPBXqGQG8
HNSW/Zqbu03bk42AXxxLWvbREm85nL9/AA5WrJNC0pL0V5YGIw9u5iJW8cyRluyF7pOj3WdsQpWi
TS6qV4sOPuRiLB1IeRloCs3oR7sfwg7SLQMdXmPGPNImks92RoaPApb+jlUVAVzqguaISATCEtj8
TIjA7NtnZlQ/ZeqJbujMOaXVSDbAfz0G3+os8S/+cncoqHCpIXps5SFXm86j0W0qM49A4IeXzDqW
lQS2GLoDeRIbeRLK0FRpL1/wqeyYNPOLm8OPvzyf2Uv2NESCprBV1f3wlliBXjfC7F2Nmb6sO0JE
rckVb9EFFsKqPC9HrSCs/J/+MAVS9lUYxlL60POC87Zsu1cnQdya7xZD5obyi7fZj6hL3wc/X4Oc
Q6pHXkPr9MjT36CwbaQj36sButgCCCXzQ7uJ3fAFj10Nm0dmcv/bZNAWQs8iOPzOzcIXCFzD9ocE
x9LAihZ9bn0clsiRCzF7h+EopyTKt6BrFwO7NP75M60NJOJzRd+DH21AoEsvnBG5RDCNHL6eheM1
oxU1nI/Fub8Mo4rTClcGCwdWGLq+NWrmUXcaVWlldKPBxIDloMmNuC5n1IwnNkLnU81RrQESjiyh
PjG6h5oa1Sr3gETgaz/Ql44E8DxuAxnu3HzCa4Dyz2z607Xz149T6LoqdgzS+Q0ne00St20+M1Zu
1+xH6Bfw4kAijkXav/KcHXwLtxw2A/DigZ4ut1agqRmHmyC7MXZIZyUQoR/p0tCI7jFbqQIj9kIi
30RnzCBczrUQSXW0nC2cEHVoyUKU7FzDme7+2bR1i1wGuLDmKe5/EPVj8sv9EkXr9jmClS3cOqnw
7HdTU+UceehUuUKQDGgSwPc8UrG5RR6KaFQ9KOTEIKOXloZltCsCNS3NXvdMZwoU/x6iwfgChS2w
5/Ww8XTEfyZ60AF4XE4iRw4oR+uk9Umsz0kTn0Orr4gAF6EMpbNUj5Tdgavy4NMV9xgVxRj4S9T8
dTEKA6/yu2ANjXYU0Jb/r3nMvZtJ9VY0r3+BI+FaAg3L8FGrZ68QeKZ3dtBl122+kVrOuBLlMobe
TfXzYJi6QTQ+C3Ao6Gel2RjKAEBIABd0kQe9dMn66Ux3apH719VdXf3PAzu+uCopUITSCklXRl4h
q0VMAf21MJjhv7XwGJ9JOPKM0IoLkb5xStYr6FFr8qkoMBMNsnLXs6vM1OmQQJQZqdjbT8itBaFx
HKzMvvIEPJ4TNyU03EQxy/S6gh14qz5FVzeE74G/4T3a0tn/nOCnABOUuBb7ClEsQ28sRg96r7G5
kkwTNszC+OyDgwIRisXT4ZxQG8+lgs7elF+Kc+mfn0feBRR8n9rKlCL9ER/rMeLTRbx/Q5r6hRkX
lU8PRLHA0I3+NVf2Sq7ZQiddTIVaG//icBBd5UlArL5zOv8oQoF8ajIhy+7J69qnubDFJV+ImJZ2
3O051pA7V+DqM8p4J7eiTCuRDoDns/EOEZTcPwfvK1zTZRPX3qRfN4o7Et1F2pLSc5VNhBFruA3I
WMPOYXU6B/SCP9S/KmbMN6vbAWYhoCutfZjRDk2NskqQv/3f5fwrorECWJrsCN+UuPodm/lc8d2M
Ly2QHNPmCuvrw9zxedif4rwQHJKQR0V70psqUD9reTEATMhQkyBHr/6tP0maLyDVviBxCJ3sKB/s
jQ3IhYYpOay7PCBD9dhf/9VVl83TdOufhNijT9ax4KHs+03pDWXkjSM8qgtbzTY0VGmVKA5iFCYB
f+0llUAxBwKX24rhPmmwbQp2DiOZQIVIX0QHr31E56V4uuFH76/5LOJyUWHiq+pCc6I9NJf+bdQx
FbHCXE048AaBtOyMDTFIKLQaAfoyLtLvIm10Nna8h8e7x9Gcjzm1Pf1u+pAUb/uD5uyJqjfYgBjG
ASmHLFGMf8FzGwLWoQsxGTyLVwsQLjxmwwEGay4hLcQZlv0e43pfwBGwO42NNpFc+T0YNa+DKcil
UYpeLKKblcREKgaMfVFpNCylaes+S39gpsuyts0J7kb0LfR21MLVJJAa6BcSt9CzqiG1wTSG9y0B
fPnC1l1OXBq/yw0gYiINQcte828PUSGp01B3uj4HkTqZzv6SdzrmvktPHUIVRgjzCHE9W9BTiM0z
E3qWzt2nQB4gPjLxjmL0o2EyR9SeWWPtNJvQers45Pg4D2QZULWVIgo1A5L3YeeZuYvAKsUfFpnr
pnP+8ND52XZIkwQndIvvsailMNduDpgSclHCQa5WR0PZg13QaWT+al0jSVF47B7MGFK2AxV+jUy5
elvZfWgc+K+qiAEyqZJ+JhCvBUVVjrxWx/e/xDQdPun5aYMYau+KQ4ipPzp7pqfurnw0XLQYxYrK
s8OOZG3jnii9RdBcOz6WxAmBLk6teEipeoRAFKUhLC0s56ghAJDJYs1ItQamtMzgTUttIuYQTXpA
0Ld8Az/RuY2YlW+dW9g4kWMS0ps4SDChQ2JoMDu5ANY65oXHIV0tl/2rF0OJmEXTi3VCHix4onuE
LCz6yHxVdy19qykOwKzzZdzSQO4uXjtaYhp/OV6udi7frRAmpbiFktFmRWBiqR1q/2ihRqm/vLJV
L7PQLgyxBMUnBz2WH6dTZCYxuCzAq7zUs2581IsdRAY4owLtaEiJY0pBykmMZAQv8BG3cPn2rpl/
PU10qZMAyV1f8kKshHnd4MAsxuv0uXks9Npcu/jF3s6ywrSoiP5A2mK/+/+XYGK7kMMvqBAAFxPh
5ktOSFW9tcdJ7MC0AJl1YRGhZ4+iSRwjSLDNdDwqYoGG6zu1G13eg4xXqe3iAX71G4o5/vXQk18o
q5R2ZlpUBQCmd8G5brBReHT3T4FBm/UWELVqGZolfMubzgwKpfuC5+93lk8tj1sdjXcOb//7jrDV
qezvaM2a7Bf5Gp2D5iEAo95XBqqDq3GcilxfnP60X60yGGp5S2qATO9yxDST46x6Y08C3KlNQGJJ
v+XImvGHTKn+yrAQ6QavZ4mQXydfDWS/7tDBGU5IuHiO2+/Rb7ogC+FmY9ABorvA7VQp7+SAIPun
+uCE5OXrg0DkWUWjpDsPppj22Yix5fkPc+NUTOguFX6N3iaBfEZQ4tmXrOk6yPHnv/IXuxMdbJAo
ciR+0saG/q8e3fTnIBMNX/3q0OzXbuQac6tCmAm++s54LvgMTu0p45LUHLPa8Yr7OI8kc4sopk6Z
2aNHvubZOHvF+OBN4VV1Mbl5a1c+ApKc07aAwVO1DLcsnRmEkgI6NSlPtnVEePJS5JoFRNan2Fu4
G6XsL+pYbHMHSArlzBIzT4GCasuonbxhp2uBOrVUIovzjcvQbwEHMMFSpZdX5+s50LkCE4llMw4p
wqDWv/u4houvQ+/bojFMBSTpxCirDwQi4R/OFAX1aTlUjp3jIfkShvrV7S0kqzE1JmqtyRaxxFAq
cTrylOxIHJe4LJd9wTdERLsgoNtb+42ENJ133+h2CeO5vWgy/VDC8Qh2JbixDvqjQ/qsjoJfXvqd
HaxEuBDYBWCUhMjifixtJ/aaDUqzoORDKgaROakEn/3wC7qHmVGcnFZm4+yaig8pABY+940LIBYl
46X2eB1jIkECtilO5QHgnCZyiiDoYRYikZfyD/1EKdrP/Q0QAJ+bU2FS6OzRAFXcumOCeKqQ1jgv
cxrSFXQnd9WPEJs3HnxB0ztqTQ1YnbJuJDh5w2tXAz/BKcHxya8TOuDEaH5IkXlxvYNi1WRRcc8u
4LyuUTqMVdXoiJ1V5YfdvWvyGMKWVtJGbb3qkNJ3PVj7QAiXqc+AAw4q5sYV9WVLFOatNfw+nXsr
qP40B4JQcCLNHBWUjF+UVp6Z+C7q/ES3jLZqOmOyFe0+I8SQxzHgEVr99mkMv4O8yxdJWIL+T0VI
84ssxTRDQ349Y7sFLDLext7W+HdznXGmF7qXSNqR4jpzODyOkflQSvqkLPClV0lRLl0VhQgzYVmw
cHP6A/Pn9ygJJf02HN8sQcqybVA2FlNqz9gtpZjw8dxXHCpAqtsISXuBaXiCADJsbTKZa0Z6FJO8
r0GzUtSOh8SBYAZiHnaYWsJJEnzbJpJL5SXGYsIGvlmjRwdDXoNpFsQnYNw+S5GSAhS4plG9TMLH
KqBEBP0D7uP4sPpQ4zjsdKf+G1augRNU5pB8NQYGL6flWh/325CySSB/8QT55D02gZvolXatFief
74gTpKBgi9+wPyVC1b6elysNc/1bBs0htxoXyxY0GeqtDYWfmhfUCilyEVTEZmZ5cU+WK0tceh2P
DgAV23JOJRNAo9iuDPXUeAnhvJIU6kYYBYyBHVqKecuGURrbn2EDmI6P+Ro/1qbJEG09xeZ9B1af
5cxHjw2e1MLeg6PcFDtvKv2hCWu/b9StiIoeInbRoanS6VqMXculr08Q309LL7hfd05Omp/LANgO
bvZFsc4y4QQSG8hryhJTLk7Yt12pTPeh7xa/AAMNpjZlY8iz8bzxeHKtF0PeK2uN8PGi2NVajtid
486borTD/hQviFIgKqMpu+NE6hIohFmGSmPVN5tNsVRz3WI53HSCM7s0ZhHy6H5QdblGkUQYeFBA
2ZQlofEuRoLFzHPyRZBDbG+KtM14NG16URascDLfmajzy9+hioTes2yTduu3ad5huuCGngMcUsLv
Zj5U/FVGqL2j5S34yZOggTNjho6QB92/OrmE03+BcfB76MDR8laFlhgx7Urs1xwCnlCAnUDVdPHH
W4INh9EBVYza1eMyQ/XoTZfLtqCn2jrISBdV2Y894WwXdcnEt7vl9LKZy1l2P1BznmKUGk9mkxjD
nrGjJCvQXJ49U/QWqWj2FQZkW2h7kLsFq/cp1HCZXiRD/IabVRCzPB+ROMEitYphCI1Xp+o/+A+2
DaqzOn/TqFfFHwgrv+yXXlo7u5e3R1h+9+ra5k93HxCgZXPeO058JU9FAz33JQRM1bZV0TPHfic7
4FzE4c6ivOfqaW19I/WZC3o+WcQdIGWju78sMmE/BOxtwQAGSBgQirVNKcskKsmf4o8Rbcsmp+Sv
NDmyt/C2ucNPKMnEKn3VL/RTBeFY52TQVkGagjILcn+Bjm8XmFDTCf/V9uJehrXDQj+jAjv2ybVq
c/VWNzbMqf+BbCMlaIWljYHDD1KaZrKU55gvOdbB4aqh9Rb9F3AiP1WekNdq5iXtZB2bxk4BEvIJ
U8e/HjcjGOQCldNmw1xFr7F0IBB+pXhPfGBASc7V45QoyQ6yRlkWe+f8apqd8TmohbzkwlGKmwdI
6Jr55qu6D8OVRFmh6MVtUR/b4y6wa/toK1iYSJTVzGdWoPG7zxpu9KAQN1OSFA3XkNMNVOdssXtV
0fpd7KQ1je7g8Anu3DJw348vVuOxUs5VCiGy6Z9LjJpxqr+xqnIbqYSyAo3fzZ6gp9T7Aed+nBQl
yc7uLN+Gzk/H5hP6pcjPPxvlKDN+RrLkR2n/H78Ld3cTc3a8kda+UkTZURLb9Sn1cVKgPqmr2N3Z
ajvWO0Zx7V4JPWcRGp742zSdrQsbUD0AOymtmAP+pfLnvc8cl08CZ8ue3Z2lb6jHSAXwKAmLVSj8
h0BQ5KVTaCXAZ/gvqvMf2VbzSxrK24VP0fznZXBnEvns0IVNt/T7vTjwvang+PpddBKLl2BO4Lui
6rnJVdkHCpqarzfeesKxGSfz3GhHnT8RFtAbd6y0J7Ih42pWgTEf0uYhH1jf3FAY8a3EjNTGBnC0
RIlCIBckKA+ZPs0+ulsCxyCHRmjlpyNFxMhWcxh9+yKGEK8vbcmLhT12uGgeEsF2zfnXfIAfeFu5
5CShWLV6H+4ru/kCfFhRs+zX+0CkZ0BBqbwhhEKJWHU+cDAfbYZq8XEz6s7l0Fn97ULMZKYQMoWG
zzjTkiYccGh8VeV2mbjkWl8Qq81vYbRgw8W1gVZ5CvWKFdwFkHhx0wpnPC/ILut9TJm6XwBmOiQn
d2iZ6PW+dWfkg8jGkA6onnOBpQMXbGzxWn/s8j4mHIize8b1VikW+7M+7sK5KHNNDi26OQnZC0WB
1atnGUXKQWcZ1FFwo8WWl+ZtfRVQ9QB+DNs48RzAEFyBUf7mfSLS7u37uwncal5Ju+rRZZBgh5sr
WHErNq4LjRUcBF+YogUOoFIc/Q03kd+QyhfYixZljByQCmeHAD+fT8k8GqZOIhxmqNPxqH1uhpbS
cpU8WQHkmE64HW+yy80eVTAlEqO5em9L+fWEhkbji2+YeZskFmdzu8lGZTw+ymGIME/my2Zu3JxF
WV3xlel3LI04EA/MBYs9aX99nW/7nKOLIbW21j8vKyUqg/5fe8tGimf7JI6eqGnAQ/hzyC/wLfWE
+v5DvsgdBBtV8aUo7Qi1PsI7bJezobKP+poDN3ZtelSLQSWQBpdImhG4M2Q1FFhgR9d/l7bdLq8E
fRfLwXAsXzIlrJ7CRe6vpjlPmKX/+6zN2h0sjCuz7Sgsp+FZjRQSBI/pQZnYZngupQKRAGAJ25ij
o7IHV7+phnHewo3uuPbqqW3IA2dLmmsrZbMBrjO5UfnEB0ohoqHcaA/bHNOPe7AmBEHbHr0sy3pm
vd+Aph8alXjGyv808XRy/yTtyjVPzn/hsOU7Nij6Cxkul92fez1T/r76syU4PpkYVyIl06lW6FEm
ZbNJENw/HyL13RnLhkKaUf2kPvJz7buuKEciBy2JhftqiS098WSZs+hFuk0ij5HczQg3xhzcf0pR
5YcH4PM+3kC7sgYsJiYTk6GgeIfVAUa3SONjKpC0FkjMsRlHHIe0kTFfs5i43/KTlImWSCPagT29
BGFv6aZxNhI/CT6VT1EZ9LnBvHWwTtu8eXmiZTF2L8GMipjOq++O2SFJC9G+74wqPTHPo9J6wVq/
LE+CkToEfZ8Y0cI1VcvpLPN8WI6KOSRy3GZBdCSrD+gBKY5RLXqFWLRUw/84kzfhiGxSiaI3IUXZ
T5rF/sqyWLMJwB30gr6Zgz9IG1AJux3ISsbKakVo3w6cYEw7u51cEYS6Iq5WHGo4nejI2wVHzoIx
a0qD1ZKl8Frkg0/d33XwuH42c2a1THk/34C2OHRoMlUfXpIAcSnkZIP2C7xBxSM22KVpbyODJwEv
VZEfLkSBXbjxGBH4SWXHKnsB0LxdCqTeuNw5tFxLf7Dv4uJJQpEsXgZJBKR/8ngisqVKqugtULob
XhI6keLvHltcodyK4GcEMruwyj0Vmz+6u0u1bkFqF75kyuWkm4EiVeUNb0lMa7yM1qEevA6OUaYT
2/Pno/N6m/EwVXltALLI7AFKrfFVZeXRyRiS0l5C3f607Q7TQLMWSlz2+bFpNlfMVMOhnzltjcbW
YotivgwIavUyErIuc/i3nkRmKD1W+u1aoDx86nfH2H2d9W6py54fZLLUUl+1hz6w9f6S1C99OmxL
CKFrhYhtPto2qLA3EeWxDpa+K2IBNadcsWvjDN1a3IMi0Ap51YYoBTZwipQKMVNCSexrs/RF9Ysl
IEApWEM+RKVu5Ri7IVUJpiFwdvP7f+jJqdeG/8gjXKoNpi0rTi8jRqUeBcrSfxJpLnGMBR3/sN1r
Cvm3QNG4rM12C6NysZ1s1hoQORKbZUqZus2SpE/ZvxdpHcEd6fwZpToG/+sTAy+LhyR+yNMbKZHe
3q6lvGUjofi0WTd4AYO5q7d3f+0EAB4HcRI391PI3FY0NPhi0lKdES2P2ZuiC0S4np+tOnEH+njT
UdfeRen6vHOSlmceicn0qy54LVWsU9Zow25CLwAfdD8EW8jXwDsRbdFjJqaIOvglHtjZfNMR/4C1
1dtHUlzgrLmw+3yiEaJHvz8sNXGlfh2QA0Xqz6bwibvKJiOVdzYjB1qkJwOVUgY/ahPQdpQy5qhI
5TRvadtVJbNIDR/Wmx8Zip6ijJtN06PGIR39HonlzwIuOf7TR0qGTPbfGNkQbdO/EoQqFccjceBr
YurCb/w+XIuut3cnJuwQZmW2oh3S9ayq8xROl0YA+X0+1uyTVq6poMlcvn5dcP4odwo+MoaOxWyR
Zd3f0JTRhjSA+AWMxjGAXicczDYv7ofvCemKLYMwALmoTulZHHSrgPhvPBU9rHvYoejo5KCfL2aY
AfhsroEtrSaQqxeO/O4xtPy9DNfLJsjh043Gctgr6ImPnijaPtDWooZ1OEGL9hY3paceQuoacZKB
ee+SZHIFXP70hsgDkMzWHP2XuHQtcokTAytA7urmW6Yr0GpqDU4H5hk8FwiR0307eUZ6btJDxY2B
fg0Cho/rslOkkAoaV1nI3QoZwYYGJvd9SwjSWrUSQyIu4sJz4j6IkxldyPk7ouxDiG4xyi2G/f+f
kcv5tEkOe8CmKPUtj6psJ9byW6uO6ZqIjGEFkSvhrfUFkV0s6PI/ChQMzbGYP/kIkTnp/vipMcck
5Fi5938mOrJCVY80woBxxP88rsjvi/Cizrk8vSjr0VGGVeqonBN60ivBRZdh1uldxyQeFUMgynZp
nuWRDq9cvBVUvzDYUDK3p/N0GrNFIJnX+3LRHgi7mxyyzCF5WAdVpL9yvAzkqtRo0qlcsr7j/vZE
fhfsXgwKXx+GtkTmnTGg1JpXf8qolvQa8dxaaZdM0xVXvhfDx/XlV2x0ij557dUtUqu77cXRg+lP
R/pcSz3NG1uZ5TjGbE2IfsT0neVLCy8g6bVw0p+i8PyCLlcjz6jLYEn9B5lYUywsVwPcmE+O36x/
dxoDhaDMgM3iSkjtby/EA0SFRmSzQlPn9AppElughw5GRN+yHS/qyzl6vwsDvZANcOuId30EMfDs
Mj8dDqQbANRKqj4XWz2an2mIj9ULiCalUFSKfCS94CubmJDnO7CKqw9X/yJwvPC6iDgx3jXFGHJM
4ESJTHa64j1bY4HA+R8gf5eQXeEXpgt4WPp8IM1NtzIHmfqEYc6gX9dEwLEknLf0QxzVdcmPpbb2
Ycay8Lw1CsYAiG2zf7xVuDLfaybyVQ4jY6rU4WFV3ewxxxPMT7Aqse2OzcI4w5mp9tKItkJkTiil
RpQVKeKt0yH0PKK4QW1WLYGCEb0F/k86W//0rr6q8awIm5M96IU1Budcx/O8j4J59dxigExXh0pj
qSrGhoik+K4Xj+OiljI2hXThqcNZtws9xH1M7cMbQQigFDeEzqNr4HuQtMWbe4xVY9wKH6dgLvTk
g2xhU0Xcp7DN2MrGURcxXOUQFA2PLkJX3gQ41wKjlWbxXKOzR1Vhx3zcK1SJXAeDKyyVwcFRQ2ko
xeYkYX5buU+LpIYPEfR/4qpBdQGIHfVSqivVBZsG3lfWBXowD/eJ2zppxfEGBPhgPTE/y/ae+A4k
Rmjs2o6WQxNtSrkFHfuF2cdoXWkTa+91AwCTH3zdWOuCvkyIlhehMaH4pAchy7QVksnvj4GEaQRF
Y77WSzLsWAdx2jEw0VG6AfdRG/fGK1TTb85M+BB5YsdByumYlyCKISzrA6IbpxQF//7VrKOLgT25
8NOjGaRr2r8YDZXCHNyix9+57zZGEYiJ0ymZFfV/rDfK35ScBUhDQtWjx+VH9M254YbP+jbG6GHx
BMSuvN83qbQVxb+Te7WNA9VFggjtSpdSnVcF/AsWD6cVesvP46BbXp/fgLrzXWR0Pew5fFoeUa22
FL5iJ71cZ4F80dG1NsEnS/bg1bHZdoofKqp2veFNc0/YfpvRhJDunBxvJbUvzwsq/lojP2I+iqXE
qAhBL+xyEKk83zrO5WAtRGP58Kk/zoU8KEa75mUYFGOxJWrBYwDu9L1zcC1pXy3DHihK3JFa5qfJ
H0ghe2bPzsJTOAdeIN0rSr4MgaP8lln8oxp8Yd0p/8FfWEsFt/BEBl6iiHN3FYbUqslhuxsGSP1v
a6b5Bco1oFunrz0LluRcpJFv4R4Sj22FOjn709bDDslSSdHtfEF23vgC4tj6tO0OMEUrDTcWfqY+
Uz/2plXWLf308xJFoHn7HlOzvo/TZFande1YSXrkD/zdBHHe5X94s106GHHpNbT2GiBXkUC7HQVT
D7k5sUfO8lmBUllzkihBTX55qIReXfzKmYMXcrLGpcnspjFgVmwXAr4LWlAb7mCUJtJj4PLfGp44
P8HzmBNjeX6/wfKwyTn9F8GbanzZOGDEEQMBuJqTKtDsjDFjUbL0dF17nLzBwG/5miikw6wkcuF6
0mZJk2cTHw5sWK+/EGJt4IWNZANWdnB/HWakdfca6zjZqAY83QEYVyK4FtVHQdvQYmQ18kkBZYQv
fN0TBz12yBdRvNmArMyZ2gY9cfeDQPZgBMt+9pzch167o/mqoFSzkfP8Ty1pTR3aejgYyoilU/Qq
oXIXdPFXSEn00tF9Iwdm95Mx7KSZPNM5FERHgxEy4ckCwtjNmpgeaxcDn237E6fIeXbNQ0TrNl7b
11ymikJzLL8Z+M9zIx2gIGONNWpTpAG4usH9UxUZFCaCWZr+YdwhncZUCOpt5f9Rci89vpcYi/D9
cfYlMjaq5+DZHRhSWW8ZeQJY4IiINex5hHgXsci/IX0vsNhqBwVHrctJX+6OXZn2l0mlCSF/AsHx
ZeeJtZ2MEbixpA50rceLRJ22ZlPDS6c2Lb3LKo9/RrC+7h9qqRIseU55WA6ohhVYK6BRrXhzot5D
oP9WOt4if29CLAdU0oWV6Fl0ms1Odkz3p+TQ3nCDbawuTR2o0ubmr+d/xymbLL1XUpH1Ed++K6Gy
BPuLUS5ZRW33ncxx1a4xGvCXSihF6cfBw2EWmK4xxa12mvP5o/40JMAy380kWLcZeKf9eqJbI+mt
FXZBIIItUwIkUFU/2Vfk4oB2n5MVzbzlB4KTuCESHyGzZgjIvjKfLxzeJQJpmAxdp7Fq8lmIUmYK
LOvpb7nNZQ82DguqfBh/DlIynpYJ6IYH7CNvBueIwgIQtWXFqXYAlkiR7M3bps/7wzZRKxofmJAN
56gRxMGHqZKmz5nK1oaMx2BUdYHAYgKpcSsyNSOg9ZVgUMVjeZRxuV/MeLHbFHQ4Kh3hfrnk5Sxj
M+fJRa0d8CkXQUALkSPtN4+PNgRpvFOALGz8RuA4meZIpk6AQiTJwYP6KqCmWJ7L+mEdoAqG0e4x
Kl8Z1VhJ2ZwPiwrYgfPETHGkMe2oUogLAZBnFWSSF9RL2OPzuMRlsVC3AAOcE9alU/1pTofeXTlp
yZVNg4r0oNa3G8wsEeN6XbZBOrhtgaEyJdjC5a7qqXl/O0EmMMvy8AQteTD3PmkNQIyYHqDRILg9
nnPDtheXCJIZpEjGNCHLwMbEW6Qd3DNoouWyMNfK+Qym99XMTorROvNKWpb4N/x5Q4wKmaKhgc1V
i1smk3Xv7KnOzEj8H7kHKlzAh7OccJh2zSghbYAOCUAwSGg2Nr3XSgPBnDQiW5K89emfwWMA/zho
dfl7K7JPZH+0Plp6YxIYv0TnpsfGRe4RvdSmHjP0CdjOGZxlz+PYLjont2wcw0D1yZwpW1Xr41Co
7Mgq6u7sJRKz0cbmxN+9CGMzY8oRtfKTQ31oQOIHqXgri0Ev6evIdQn5ehMZtlOVbVNxH5siBXC6
LDqSaJxXBgkbhs6pQsnzoKlgbfG5dSQcvueH4FWaZ+IhrXov+lxZR0bWlLOoVoJqtE5f6Wp5Ofev
9JjIJZA1QjnSie7D3TmMIRIqKbttZUbj5z/rbqHIXqGspoqAgj9jpQcD5iODTgk12X3wIkAzwKof
eRUs6AElJHCiwWKsS2YBwtK3PbPRj3h5IQEaLPRpOGm+L0/tE7GgONjeUGLAHrnkTo4huba+O4BC
MdETlVsVYQ4A1icPnX52Y7CTOukm4KodATe2EVqHbXZ9cAmxa+RBZ+a0wGEmpkGHjNr0b1L/4vR0
75ttxc3F1I3diHcSmhW9UaQAkCjddX5ef9WoAy/Ev+VABvJSH/Xrrf2UeR+S3aEwx5lS9uTyV06d
el1QMjdRKsRD+8CKWGrmuFu87JsviZ0vGXXQbH3rgVwf29uRhQeUPn3behceIKBwDJIMfOWna7e5
3mVSCZZs3GvS1K+5Rm586csuJJXcpWhbMn/eWwDhCASfr+lpUp6oAnA47VlaFxChGw141iHduf2U
wVkuyBsdqgOZf3CQWttXtUUN3cdMjIS80IFlzhCmV1URJnzIC+dQ9ZVCQkFHktJhn/fna+AwUbz0
0hA7XLId1pppHgSlbdBYzGBiHZJAk87tiO+nM/qGVH/4dpUxj1UhXNCt+CzhskTgqGqjgLwRUOvJ
FdRMgV4w0kLzXOPBEu8hzIvwRGs6EG03A2im163SZCc9iU1mwIfko6gXiadWcuE+xWDQPZLhs5lJ
QdM3gC9AoL7eoE7MdkjhbLdYbFpvd863SgsRGgi2Iwl7j2Dl9ZwIUjFlRrcaj+b/baNXh85mt/HE
er1mE1fcmmK6LPySCHjhAUCTClOrHQAHuDazbwR91cmCIYOqpP+90Ohl8k2DSi2gHx+CjerPxmJc
S1Gum8QTVEvqufJRP1gwJLNolDBdN13oVgKSrjlfwgnXWrk0VKEw3kOjtoGn8kJPkXVwpoIVXYCX
9ANKOujbTiOT3SVZhJtjUj46lMsPQs8LfZ2UgZPIy6sQ6DFFglv0kEIFL1u7Z0yHAYPvZrEQCEh7
oa3/TbVJ4HRxjrDYQEiIz9BDFjfFQ6L5gw4eUEJK4FQ+7HpwEOSUPGdU3us9NDpiulYnyUNHZ5RD
CkIHYwqzv/6nZOJ6Q8cFtqTU3zGRAYoVrhzQZyEiOnajedtQBzkkvmPx9v0xuoGmTfz095nRnpPU
fHivKHwQDpbpGDYu/0uMG6ZTBSYDFesaloBVE+26w5xs+phVQx/fe3uFBVUm4BwV6qrXF5D3Y6i+
wKPuLARA85iKC1AqFzEVS/S8PLhvi26SFI+YKSsgbhemQ4ja7IyizPYQT98GFXhJTzrL4MAQsaVK
Ys2Q3Zaz39BoIiwSQ3viujSWFyHUHVqnoz0KAQKrRqTIKSgIZR9c0/pm/zHAp4Eo4+e58RxmkGAb
TSyOmZQ3CXBK0YfIk+BAEMpZg4ZoAG9vIR2lfzZbCCb7CSJW+kJNHys5vQYigEXbguuZeTgE8y3J
aZhP6HmK5NNjVwT2hKBTMwf14qKBJgx8vP3HGOhwdxufKoiigAz79aQFfl6ppFTNtkh47FUpkpdu
obRI9ILx9ApOJ/ItTdcfnBkL562tMpclSgn3aFjVNd4yA8sHxjYlinq59ZhDmSoseFlClOtXVpOU
yiyxpwStOcSinEOjKSYkTFc1isMHXn3Rqjw0nnbkDuuP5sb/y3oa3b3qYDBH/D8UGg+001nU9Goz
yU/ghGtfZjtD5iCTeajSxRPTnlm/iH0zfKYsxRQ6XrMJj7P2OVqVNsYU6uqrkDf3ZuYrTHnigWsY
vlXEoFkI3yk2j70wF4r32deiOhCuOXd+haOtKqfo4phs1QFSPy1OUnoofXY5MzzhTbEzQKpnyeiO
Wk4bhzB65ybxKJwCZDXvWZBtF1xkUh2pid6dL3jbxYS7M/QSrfCSgZqLWiJ0k8L2BL9cnbsWszl/
m3DzoI8JfpDCT/6CAbR9jGCwG1fQYfNsNNMnVM2VUwC3b4QDgNwHyh2a8KvypJIU7frKU8QBrxlj
wHg5MwI7zFQ741T4J90hnTBnqfGUkUi7QdkHAZUs4KiaDCKGBJoFnOrOMEfKFVF2bgEfxVU8eZp/
gV7rZY6CMfttexlTmnMeKRc7dUAKoRyVM2M5IuND5A521WnoPa77PVVk8Prv7EOA1+4scTO6IU4b
I7y46eBMTyhDVassCgiu0JYUOXNH+9ON4dVlB41EWgktKw5a09V5IB6U0KV9l9x15iEhfKyARSKl
m81H4D8ur/fjXUEekubxWT/hCexGVI+jF01LVeA3VBXedzeLLcEeE0AKPOgyZSVfho0WWo2chwmI
RX+aq7on3R+9umAP2TutRoBpTluZ94Vv4NMdw/wWWg0lHQTFGOWaUa+SxLbjZgYksk7rqQxYiuyC
1NsEihUOgEkcv6VgqWAGhN5OIeTDgBiEpg5+vwRQF8oy8ecEwJ6iDyyKiyzjqa7LX9tltkAKMcp9
zO3RFc8ggSbtwnn2v/EEUTCPFByHJLu89nZKYHlYvzWGIMr43vOkcsextRpgf9/RdIN9oMtIvaJG
PpbGyE7MYxjyH4UpeWmrRoz76rOxqhBC4OR3BIvt0Ndkxkiaa24IJu2rigIFjrrditMeZHsuZbYy
eHD3T68VT6qohRjs754E9uayrmejr4FFHdhHvX4L9pU1JcPziOoejyqbfUYS/ivib1DUZ3uz/u5S
jxvTs3Nzmz/cjRf59PUrdnQ1l5/2uQ1Z/8ehHu2yZih/nYGVSs/fteNp4OWSjqe8KZgrQ5kmSbXn
+KqOa4bivsSjHCTN2Qv4cC7uUtsbb1AaqzRIBQS+0bmDbGwzpMKnaClH5+Q0RMWFYSn/Z9orxAI2
+6cAAMs3raVfbgO3ntlHn8dT8RqJHai+YvfQ54VXb3KAMvir7/a38tjrno5j/xBt2OqGTRVFGaIg
vxzdzQNd52RNaAdnJlKijW3izanmxtfdBQMxACu+7fw0DUT/lKwp3cojw9PD77vV3eYx5DrTIwjm
jzQrlPviMQm0OZZRoPxZ983gEGE8aVpBqUMSAWIJLj7bmuvRv52W5FmZ4hHv90gVEJ5nF+aygjqU
oEGPEsOJNqIt39lG6h262QSKu6cTHDfvtUeBp+XSNPMbHQtcwnVJ6td9vCw0rEWRcg6zhEW6wx/0
iCDUIfNydb9uKCw2SgUfviSQ/wZvFTxDWQM2Ar4L54BKCSSSr2NnwfrLbeoGvWRoaPnye0WzyT2R
Ao/o7zz4z0WpHW/qgDHNmX70x93ttsn94RbJXpCpnw/9aDCu9o1S5sle95cY7eCy0ItcGgQXLm9S
USZ9QlcSx8dvhdI1q7Wmmm0gAAJxvkosSVqEJg+r5SToS2kA8sdTszLt/KLI6W7+3EjSqdxzyuu8
1t/u923fxXQylSuIMY/9Oj82fC9dgCFeA1gVzJeQnlKkt+RirajpmWE0wD75FuSFB+CPQIBwH8Hj
a5KL4ATI/CeLyl+Shlm7QXDNmrQFMklpEKKU3Cl/gWe8q0Y56x3loxEfrvLtPtKeTR7rbrLrfFVH
/L4V5vsINLOkPdj/M/HNDV5fNlUu5j7nF6hxmN7sI1KuJvXJm4ivngaWeed14jr7FUVeliWW7BD9
K3pI5acLoIs1siX9F0+qUb5wlohyxGGwoTw/snVxKQ3bhpW+DuCl160fgwiNT/a4/FiI/XoH+8ov
WlrAOv96+R/DUS4xjpu9lIWWaZJZ1Tuh8BKrqmMhCmWMtPf3Ucc5aTeDXdYKac5ZjO5TLUJ4ivaT
N6qJsV7hhyo8XHYC0Po/TI8DPRIJn2b7QVETEjH3Ir9W8ALXAyjNLJC/i39ZdB9ZLU3m11YStSKR
7mirPLCMdPKkC3NjVeXubgutp+sDvDBJn2hrlU49HvQ12DYMFOJudZFC2TI8rT1o7XEtllPY8aDA
2Kx1LJQWttT6HsaquZ8dzWO404EBa3Sdu8smUl9iXuBr2N4JZVt3ZEJzL0cUawVuZDYnFC+oO5IO
uvF6qoKF0Vxki2B+Z8STSwtqgw/yOH8RwhPHhGkOz6G6wJdhD46kLPYiBKmfgLydNLNykxPfQ50J
wageFAP2cX8oGaMX9ZZBtR0xrqPkXW/fEq04cDXvHfx0/MQcNaAnYTZpwGKpmSSO4RUNZeRYTcC/
D679niP1014YbB0ib23JrKpalHbfNfUTBNz/nKMtp9p5EE2jjRmCD+4d0hhifwh8iix5F1EYrbig
t6xC93+UV3UdcLM6Sb0ZV4TKCd5yBbBGHZMuX2R0ibEO4yhP2omowmLVMqZbbnBMnFLlXFUZfqwM
LVUnFZjceAFJCL5CzVfASnOH1oGYpqDgsu0jq/adaAGzo0Ix1WZqse3Xe9GL3fS1qUXoukMwC8Nw
Y8IBVz9b8+zHAIdvKSOR7T1q1c4gdmojHT1RdinFA8vufn3LsaeFveFUhAulNwAGv4hfxZu75m1Z
Y03HaETNMLFR9CIqfAxgjBIjl3UCVh5dM4X8WZhUB2zC99leLKPio9QGdQs6SN6SrAai3Ak6Xp12
56RXQNgcEQAqg/ST6AmQPkF89qauUG8shuEEJIEYB+TzIj1LT5vYFGHqVPYmt/gQl0IMOe9UFn3N
KflZizmsIPnuXLS+HK5XAo7luPplwgPYQglnq8DuOSeSeKmrph5RLv2BW/Iw8EH3oEO6SYwh6ZqE
/F4xUciNVza2JfByDzx/ZumCIyB6NscZxViMAx/tOmO/A/0z9ahnEmaMrPZhpcqdC+Owm/NYZOZy
TvvYs/leQpk6rPv/L/OJ84mivoZCf9fjpADYqdV/ACXOS5WLiLEpNGl49IlixTeUTbkqq16PAGSi
zc0vwgEDZaqN04pjTVcehER9u9MwMjD596Gr28f0Q+zJagSoc9tfJKRBj0r7PKBYMoQm1EraTPL3
lSN1dtZoazYU9mGDOfiDJqxiz+5I3xmeEjbZhsPRag+ZPjn31L2O/qPmDY7P/zOPqJIw3FkbXxxZ
KUpt+9tw0ITdTGFGO19ikEZ4Xf9VOv6ZaxsW8ZxddwtBP52WS3zQBM8glFQzTsY+iGw3HZLZBtUb
JC1MPrUD3x3XQJ3U+He2b7FGQjEn2qMqktIVw8r9GyWWXyB5raTzxxLW8Lqrk2PxquyJAxkxuPEo
YgR80q5X1TYU6luydA03sA1fH5HqJTdpK8wLRuIA/5EQ2yomLOGXBtmrRTxxxECK8t95GdSkgmhV
fYR2lyiO1EW0gUGmpMSHhgLtvozeKz8qc9wI8RvKzwoTrXKUbduHVaKMiH690FnZBwqmvCO9eFVa
jHte84QzDxkL7PLw9O/t0dErGXtyowZOwny62eMjfXgXbrQXQyr84UfaYwgBrohnSSug/mVUsRjT
jQ6g4IecMqe0ZaGvapOFb9jGI8xaO+qaeIwMAykTUrA765btytZqwno2Is28uUZP9BqeKH0C64Ct
Qxox01BRPEliDK3uK0ZYmW8RzNngnzKUefx1ZqBbSFkGK1Yu0uEwiUsWhA5CUocZens+pv/fe1cx
xylhDGgKr0qMerKlF/OF6pg0JMC8VnnERTVVolCN8FCMqa1dRrYjcI1CvDT5XCXcysM+deGgHOh0
Q0P4+EiWVX2y1xHrjXQIFFCy/j6oZsq3vA7SxyD1DT23HaXdp55ZL7ZK7+NeDnILi05hcnZPT1QR
iBFAVcBuwWwALFjKmm8RAg0a8pokwK8awMwE6KnD8FE58mW6fdF7A5ym6iW5Ao2r2cOlASMO88FO
rtisTwOAfNXcxmAuxGfR/PgBygx9MTi5YYeBoNJvfS2wMUmuvcDYKfhbAX4+hwF18dJO2AdSc7zF
yTjHysnxGLUkGN96KmyKkTX+iQAhy6Mi77kA4Ds8oyD90Fwdz5aNi2VHsaP8b13eLIY3qkmGK2TE
nqAF0DEvK85MTdX8seRYaHjN/8HH4PiYegoW6j7sD9eP9jQ7M6TgqGV/3R6x6l2EtPU4tTtlCkU2
AQAlttcJKcZDNdhu+T8KgPE3YZpEYBB0mWF5ZBIKB9xL2BT7FniPxoq9BcgX23Cn/gTmhBTQ42Ul
aJVjbxvUGFWlmA5PtQDfPOv/ZrVYDTA8U8Wo4B/u/FYW6zDyOUqiNV8qigR+Zn70ogl14nprWL4N
LTh/Z8nGVSGRXpvijYIECac4M4OXjSN7z6mR0fcZPW3RYaimJKBc7NmaEw3khJh/+ChsXkZSi0Kh
Av8936EQoDdzez9cWnXbC2m7EZOSIr3QTXXE/wySVWYsEEHq0LSmFhlEopu3LA8SM8gDRecTLiRL
Cv25E3RwgGdLg4Gd0+JCsUZxGADxiQeerlwy6Z5fko1RXpf5/ueX98PWlz+3OE3Isro5s95kuLNv
JXvJVFmuVWX5ZqOtuNLvin6NbHe+aEuPGhptPwAUY2W3tOIZGWVqhPdqPluN/nJktXVINOcspu7n
Drj8oufdr9fkZ816uTv/iapA0VDF18i2poXvpPELATq52GtS1QKzwbhQwrtIoNahAz0F+El7BaQA
GZZNPP/xxX57vCHLeo74sl3h7cnHnUPA2dqv2jHVE3riq2GlDbCe8APp3y7GpTQ1Yl/fgsT4LLGS
qmReJVCAjxDSt7Tgfo5KpexVGu0C03k/ph5m8jQYSRvubOc4VCEHS1BUg89rD4kmKc9TxCqwng7V
6Yi/wVmk+eHFohHXnbIsUcmiDeB40n1DSaWm2NZTJJwxyJgsNIc3cuasfBtF0S0Gz+72cCIFTIdR
etbA4e44X/pIPa2MPRMrTf+Plk11argF6TZpsvRFmb4d5auDGD0KS14Yt8QarjUaJsyuE5Ze/9uD
kPVZCpKPjTkIztsFGk4HSxAB53lDF3jhDT6hyuhDjBleslfvHIvfE0sAujOR5NF/P+CPJUSkSl/Y
Cxq+Okx3iGPFGB5sGX8TnLcR+vm9caTuWaAt89SlhHKXBp+ojs1IkLP6GVxdwIFPEqHDKXnY4MN0
0qOdYRzWb4N23PNoitnoVF2Ngk34ctqLJ+pE7uXB22gM7kl87byKt2bS73Dp9aAzedSmunyle1ym
OCAG9xZ9r4NG1xrGLX367HYbRaC1Z/cqyt+aQ/g5eH5q4CjAhKIBmDMph8M0vNivHmZjSrpEQ4zA
pu2hiGfvNIEoU+863fKiVER2tomxkYItZbk/wQc2etnE4nF5MNR0DmVkyrmwSVHmPKDptL2VtHdc
HwvQzXnmWp+fyuafiCbGggpar3tI3i7UZOJcEhYOXTzqXITixEoSAc1CD1NGTE5uFA90ws7OjST6
TtQvohSylTgIbL5BT3tuBSM7UnGTMD7dl2xvijb6dfufhfP0nH3w5JCIprWT7uGLAeGMyOkJ4t+w
RpybrsCN33dgrx1TRFAXlHefZQDpOiAp+qArNDmLxr1TC6woFc7TFtTGGueN+PSG29s5Y5TOZLMi
Co5C+jQPmqzEzNVf4s1hxqIvqKu+579qeeIU/QbrQk5X9Fy1koiwfkZ+cPU4zrSMknj11KkAhrvO
2hzgE20V8EJVx48Gk2k5yJ0FKKq9bAYZ2VkCSTayqcvChcHfjte3k54el2juKoho1Ptw2sKadP6w
YOSvG3FP/BGqokZA6tT2BhasxQQ5ss/npOqWBqLWehjAlfXjRbNI79KQB92q655BowlakqJTjKI7
hONnKL5xIq/px1QXjbzKo/GAADRlpurwevfLs87v9ejW/HxmNQB86H8f7qrXpkLQpCvfA6TMpzMo
nn71K+Q66AIW31bZ+tZELikd9wxgyzUGt3zhydtsYg6sZFHTcVPdgNtF4d4GjmoGqGadrJtVLX2w
1xSJyo5knJax0QwdkccVtsUhkbesWKz+7tjgX/dIBq+/cnPiXdldZpOuSkRPQtVOaK3TxRKeFLSq
jvkJGtcFMLMl0uVRKN/pbGbRvo5WokIfu3DzXAGXe3mcOWMvC0g5ib2+5wuB7kcnP65lV7tmtrrZ
9wyCGVPHKTGqDlmtOnElaqdCR9FI7Z9RQ+SYeGcSF5lDPFLvWHqBVijQm+7PKdqxgOMprGjIdIwu
NsogD+w6amVSpT7TbYQQ2iae7qpdLez0n9uZYjx+Bjtt/p6pdIPiU9FK0vEBeAsGOlmf82KXcThZ
IEi2lwJEEhuoq4PEUcdYnBAH0OLFoma2bl4NqJXjhscBODj8efoZi6ngt0NBo1VcbPvP9HWnc1kx
k7j7ThLbjxOg68ZGKEVb6Ax5dut1KyoOHWGns0VnX7B4nQ+KW0pcTh1WNG/y29sKJ7G2QjuHBL5S
ZyzQycaRpx7Q4AjuFoDlCi7od/OOWE2udUveEkzPazTY+lR3wJYYOxTxAnCe0ESllXD72B5CeWm2
jaxxrZSN2zRoL9uEpphsYDlMXKiY9hVYZBlMee2UmAwC8ciCn1Ooo4YmIRbQ/OOy9ZA9o0GPoMED
MmKzedlXybz+gSBJNVHeCrjMgTlJgkq71ene2YDAtLk7Ov3fkU2UIWqdQfgSHlqF5NgY+yteuPmU
qkl8hKRbCKrPBJO5cU8MNxT70Z0O0oB5VcZlsaI/grS6dZ5F1VBe+qrmIcWZJYNNXs2vDRp74/AP
P0wnyNOx5+3FyDmKQK7STi07F/nQ8kvM2nJszbIeSwTm6ZFbQhPPIjvz2rkdBS9m7kvyVv6O39pn
odPOPepjiiukTYNPzjLSkHMtozvpWdEfZMfw7NG7EunqJvuVUF7jBiLTgZl+hNZOZW2AMhMfDluv
ongZPwHGECegdJ1dBGjyFuzS9XdBRjVrZoVEU8RDoLBm41NcDGRIC4PKPMVtTC71AR/Dn+Cb/FSy
16UQVRV34eJMtvQiPoom+ni04qob/vV+LesPuqcdPXlL5QGvNwVKejz6f4IKX0NMHXCHkanVux0Y
Fe+RwQnAje8YHzikFmuvz4mTjJ2pjYF3rKfbDZ1UKzMaYWQ80qwErHhLvNrDKHTi9rmDKnAThfrd
udQlAsE9CYonGuT+SetZvr8llmAXUyqVBKejRJsLSRbAIIXdBv0sCTDbo05gBOgZvkxDzSTW1Hjh
/TQHYHXCUosbxDBc6bp3eVti4AjyVjR00SlTkTaQzo/RJWQBfRAdHEf+qSBad+h9LVRk/1iJtq1k
pCp0s969smfj6f+pU6KY/i1XE6rXtanBmbJDBGO6KF3qfbrtxaBV7LsHR/hWV70LMwWlrl2Y/IAZ
IBB+WGKMY308JUOT8GgqDw6sPBtQnaZv9y+0+vOFHrBqntfWl92v6+ys3oY6+7SdOAkJSvXVZJbr
A5Jz/NXBUIfrccaXOwyViPecPzIaChccmNd7DM/CCYHZIFbxpp1jnY2j7DQbg26UPoaZIJT/OUQb
nONhk6KjGdcvSqy4agBmQ5Vapid05iPuS4zGSIZDKm4nQVALWwIJeobNipc7KWDuVCGJA0Y4tTCR
+Po1/Kw9MtGlgBxo0HUDHgP3Q+Cl4UGfPkMirYubTno6bpoUSfzsiiRjyqTKOQWX1cIvJDMDzmdX
i8PYhgfPxcV2NQuH9qjc0sS/fB95b1nj7f+My34aDhhwZp+F4SqUptqHtYrjuraxlhgIKs2gEsGI
fBnOWnR8iqS3ZdSQarV2vRptFfyRQTDGVZJbffRJ32mj/joYYaf7J/4tuvkYK7j4Gtqr74J2akvr
QohsLMvfFa++Tar9lfehkcTDJmEI6NyaXAgag2HyPM1jNNikOyOnHQdnRymRysxOlEpiRAHxCfvj
J+c2289nRyPqaeC2EcVA/AJfzVn1udXBypxys4FmETvouMXGVhnF2o0vKvzeKqrbLRny+I6yhP68
T8mP4thkGsT0jbMUj2d/CP8kNKgz3ol/85QLyMAXapwG4erR0ag1dIkjUc2EHGiPIMpqSFGSAKfm
/9kZeiw4NVKiHD3xZFJcknKcg3UM8OSVoZGRez/nFVGHEL+IbTsefJFmDcHWmZO6UfdeoNyn/nGd
veZDotFTmFVaov8zsgNZdbO7c09NcK/fKCs2FSSeQRPpVu+gbv1XCb4JP8sMRZA2BR1MTtfdlDVb
Vn+ljP1h/t4PJJUgaMoKaiNvcxOCefLLdmH63znjr3Z9tnIUABEtvsHi/QSdvueYzYnUktktPsBY
pjU+sVh+JcFl71JrDBZ/FU6jFtkq9m45/fr4aa5zrs4jpueT1UalkoOaZeydc/s179hys4d/aAIW
noExGhe/3c3ioYrobMIwjdOVjvMPCeqhDoRJqzDT6ElrzJbzOgG3roN5I3y7GSBOFRvY+8o+EB4O
EZdZjkcTqAk79oNvLM1HFeAfHJQ/34FSuE6ohmH3uYdxxJ5hDqjekmEBb/nvtN4192C+m5aI3P3Q
ZG5nfhJVdleb3zFXAEq5diJ/lK76Li+0OIOep8i4pgG12YKvLpYSxQokNUEkLUeZB9LznnrnwlU7
HqJ8qe4ii+ug+dD70Wl1bXQ6h5vfaFE70TXUmDcK5xR+bXj0DTjxgZONK5FKB+4St6HqhiU8/Ii9
Oh9V9ZJIFbMPdqmzB+Te5g6CzggQf5xxj6PJstq+/Sy8KZtesJtKRopw5jiwf0o74QuUh4z8UIuQ
awpkfpzBZBgn6rm2gYlQFY21VsnRg1bBDGZmRezxsJ2hyY+xUoGWiNHYQVRSc5KwurNMzOULhc71
J2plP9Bi6/6LCknVFo0HM8QTBzyZkd8l5ycOxxOLJNOB3cT2dCOq7WqTHlpppsOpAghsjpUBbJdk
Q2NBxvTpHK9ORDRTX1qzMk8VcXy7NmUZNEwudm6uMKIxh4uoEeWoAkzrC68fgqdXC81Z4NWffDzz
dBDMQkuQNBSjMSy+VTi1bL/u9BNmVg67KxKcFy+iUK3WnTz3xz/OzyVZF7OZSiHbEaIuAZmewlTa
Id/vXE/4Mtgv8lsbOzUsEYc6mLXiJ0Ba1fvEurJT/EAlBEVzgaidTvWQ2K608zitrRUp8VbKPrSI
0/OnpRH9ZqxKdsiLxIb3P6/JqPRVZ79hrWCwzokAUyBx0do7sEHpGx1/0vdSQf3/4jLpU9xCDXSV
yNUcY119FL+JrdiuImY4kfk7E6nXlvEPOmqyIbpFFyJC0sYmfdEVX1mvSfA1l/jsELpao5wvEZJv
1zrVaqzFG2gjTbXw4LLpedEMuYapPmkkTX4oRW12hIS9n6nRtud+zWFoChZrGTCPX4/eh1dLCVG1
RKr8VVIJWcgGEk2z4oQ0r6rYIDr2nmXrp58wHDX+BAr4T5Ly17/NHbBDN1C3FS1pL/bAYRa4KT1O
rgcGitqUFxlBTWhWTV96Ysp8XGZaJGGRe/ul5aBiWjWUW/341i5xGbS0SW6u5rdNVml1crXiABQq
psj6IuHpjV8/wAXPsDvyUn0V1gakgOlsc66sNfSNVeAElHNA85HcSWX9dO7pKCPWHmZ8B0DuPnW+
Hl/9HYrZWPGOl/vufkEOkdwl5teAZRocgQlgy4AWkD5e7/OzjzsFLA0fELc8slmUbIroQAz+ixHP
9OBKGGOZut8m5qr8qtmvofe2Rp143rbicXmbn9HBeRBy5aIz6/v4YwuxMQk5J+KYA1Vtr8Q8yRCE
lt4oD7BJaO2j5LLPtN8jJfidBHQ1LUUaVKMSRaJm3LsD5151bXzgKbOcbtJCQnB0rmpUeHhrfklL
+0Dc2FKe9dDQRSrSFwoRZO67RH1r7kZtshErMcOZYh5BJzPGSmQZkkkUNfNdrYsv6hAufOZg3+pO
g0SNFtA88RCl2ay+nRNoToAPX/onIifBIb4mql/ndAX3KjfafsiQHmwOIXHVpedrdc8RKQ1U0hvq
/wOAZwYOk/mwFNaG9xCRAuQT7O0h2xEHwlwOkONpMZbsJ2rVrPU9G3dfOEMPrUk9y/MolRpddvCF
brZ84xPHzmKHpP8nT2E4ceZZ0798TA9hXCo5rffO9VmXItgFGTQbWKh3OEj7egvwsDmw0HCMmRmE
7fbNsy+dPa+oxXcXuatMmMYjnY74mZI8ImgmQOcORQm2tG/QjkZj7AgJ/2xJHxyBj3nUlBo711fG
NBNdNgxAR2uDIAD03wG/MlCCQCR5/frD94gM1SIN1EW5KmCU5Nh0Yd2d/W7crXAahH/H26TGU4Pi
pCqEs4XIv/zjU6hf7gliZ2v4g8WBdwFxnAVjeNEq0N4vZUCAAh8klcrU4EYyBBBkB8fZvXqWZ2Ib
mtu0xhbWTy3K4JenTuq09rykumuC7wAuNDYSnGFZbHzSnnsaEh7ViW7cQuhtQmR4XKXihuFWipJ6
X8F3uP9lv060+BfJw/29McYCIimq3URdj1onz3gnj8pqITJKo6kmIHUdKM22Rqw0dXiNEUyNAIzg
DPCdH1/R2wdhJYBsE0/CADAjU+oMlLnSMhENLBVMt4DqGdhzPx8hMdkKK4Blq07v1Pk431+QT+Ip
VkV4ydi9kV1P7EFzP8jgc7xCBT4iIQYwBjynHS0v6EcNLCTjTM7KoeSDarCP2zrXrmPsW4+TfdNB
PZcKLg7fZsPsn+1rT3mY2azsyneehba3vPrZUXrE1KQo4nkzxQGundYG+7c1571Y7WYHWFcd64Cm
rX3gTUWPyIFadhbKj8U9LF4hFHKd34E0OqNyGAOXw55pmgpBYhA7N+WRb69BplosnErmrlna4ArE
McsdQExt6OF5LrTS/IgDxbUUCC2WTUJ9/rZnT4pEGcA6ZwUG8Kx9pGprWXnIAj1fMz+ys13+yZrX
VPXSw6kcmq0zbaMKxFmZ9LHGdN3LsRkw5UAymcG61JRjBXQZyrg4MqBZgEjGmORQjermOeukGFYY
4mc4tOHaIBjm5/Pk4wcPwGGMNlrDwtwixMu4+D6A7wJOiEQ+M20QNFJbCyZx8TLJhhwTJSrcDyoC
5wKLhYyHnyVhGHUgSoKCjhMnqrggHx9NUEwneyoeY/+XHfflFEwuzdeMzltliXSx9RnBwFaXpwU0
rX0JkbpUWumKMK+GZVHRPQLb4VWg7x/4ygE489TBhChdoTFN1b5TlVJlx41R8QdFS0YzmkahhmET
+itVukldtOny8x4rw0a37r5VyXzIZJOsnsECpRJSSf8BFLwg5+w8IrzXiAfah92qyv5ehg5Kf824
tRZtNQiX9BmllVrpm5bhbZTzEjh42CGgCROn7N2rkLeORS0Vaw3y2Y2QFTUDNdRLW7W1n24M15Lb
U+cXqwhNWnWo91sYJ0Qn54sx13kZa4CleonIESuzYxa2goM2XIULARngCXV0yfgDYfuVyi6e++Lt
Q/ezdzNHkmbegCkQKgfWy7Wsu6FHXO5Fw2Yn9Lp3t4auYOmT2nyrVDsfngug+IOH1nxiU3GWRE3F
LhA+n/IXQHASRfWV2svD/RyRqneW6XykC1aIn9odetH5knbpo88be6nlHuHC3Mp/gHn197z8ZPvV
HhA+ROcLk8todA/yF1vR1F1YWNHMaDjX5yJQ5IDHw9iS4+Gakpw192i5l09gIvsVEEsHLoBPfiKy
WX5VckxFQf/uEpDuCd9vUnQ8ERPuOgdHH31/KLS6ZCiNHWtcCxwQMZoTTkfkJMRaz0OtxXVegmys
WoEqRLStW/IAPPNwX/AwvoZm9dHN34rDO+6rfEkt//B3EjPYyFDLShv5bKuXyutSJPkN0M94j6Ka
VfGaBGFx1Vk0C1zFrKaNF6tWKbwYBVb9gADrwl3LM7wG/HEHWUicsk2haiIUAumQHzfHUDg61ppa
bNqNCGikGxs8W2cYSBfJTg4WIhcvIw4fO5hpQZBreRsdLHOiVpavMJThA//So9PM9k8SxqSJY+Lp
STL8KLce8Ke1l03oWn+8rRtyCSRfqjB1nix8TKENoKE0YaBMSWEDM9SIlivgAt6kz80cxTT9/P8P
PLP+10GFaoZ5GV7LS/uJax+1+HVdLF8L3ubM3RVGtjR4WD6WBln8aD/AiPPSN/QflpkPJaAlNQFX
3wo1ZUD5vwoa39GGJaDlLVrVMJk8gLxHBvUqcvPNIArlyhOC6T2oM2YrO/1fgyUBccZsZ3loIDEf
EqlkZxjGMY+9K1JUEA1ku8LgUlb5UiuggDcvD4fVVsukEIM0VhW2ANsrvlvVBWmd/pCRm91wiyBa
PhOjstMfyRmLycQ9kUP1dXgcRQFXd7BfqoWjJLXwXKIac7KS6LLfp+jl9Kci4V6P24ve3IUSf9ft
iP5wIDCvxXly6+RdsPdVnMB4Stubi1gZhfcEnRi7Uud5u6Io7522PF5VoYagJ+GNrKpkwA/pNbzJ
yKIfbZSSx5yITzYQydbWbN9Bu81EFFAjcA9178ZMDl4Xk57MrDiQtN7U4adviOqEyCZatL0j8uM+
eDDdtGIND8a3H7EVlRrhrpZ7w+EiDcykhGnj6JQi2ZM9AAYHNShiV/q7nJEm6lJkGFAKk3MH6JqO
9HQ28+Rj6tOgIwSF0EujiqCia1+sdxH8WbWSN1HiEGwNrMatqE45+C4h+QeXecLYJYpIx9m54zc8
5gJ8dGOTAzKRhuCxaSckNdHorQPnvxpMNS4MukkOIgjyOqR82UvuCKTaEfz4vblkc52BF1XWrZaH
87GlgzKWlS8XMVJFtIVZSA5K32aaTmQ8LUIodGHaSLxh01MJO9W7lhrcuZt78y5y3Ectm9Ay+7sT
4clwFf97SQIOWwK6jyV8o+5npnIAKrIBtMEzrZEVduTFTsg776uHUpUrwAkdtezPj1+JsI96iSTJ
0BIITT5uG4/6GCe7Kp7kl7CJFG0eE1XkUES9ugN6BcUssX0h3obt4VS5GRyGVIswyn5NNMavGv7H
LdsNvBMNcuL15dyTIYwGQwRfTri7sjyeHqeAY47p9A3dI6S/mdxfaff8iT8KrEzMHardZQgGKqDI
ZYoleU+hdAB1oWAko5CLvJBnNAmBmJFBJv8JNnBWQdrLuPOptk3iJ4BiOFKP60c6JKi2YorPn1sR
MTXecGrQo/gU81KFYLatr37pZsDRl3nGCLBbQJvbxqEwrBTO+gE2wUlRF2DBwBu7u7VzBZNpNUtM
FJQ742Zy+ElRgzjEP/4iRbUaaF/o6Qh6Rtp0NQL2WVfUrhdGHZef1WH1lSzEpLxECuqDSBrT+QSQ
aoPwM2w5P6tkoqkszUa5nJPJIdo5D5n3YQZYN4EWxp2W0zj5p6H7ZlWyLrY/hvUojUXTX3k36eke
m1yXlrePD+sf006Pe0obCifm5WygQn4WLn3ebBtxz4MZNI+LEdRK8WkOdEhs9Kkx02e9HViuUgIa
i+E7ZIlVJNg01EjhcrO8brCMlgAUKMZr37ZcN1dqQhZvL2Hh3D1kwNj6BFg/IxarUfAQrrzgUuQl
qoiRNqKSn+IwC0ndLtEOe9DcAfdQxnlMIcasYC13TBoz/23ZhFQMEyu8VaDCMd+DoRscTvu3gPD2
u9F6UEooCzoqJEvX7q7MIK+iikyLBYR6GThODZQTqF33pQu9Kveb6RdsigcVJSxQug4bRQ+E5Q4F
aYOlmd1cLStHLm/0YTK0G9d+H7wmLqPx1gPeRRVUyP3FWby+KXx5c3EfdbxLBQrenha7Wb5lY3eO
ET7Ounjx80TsjPR1O58sXCni2cDgckJ+gZJumYaw+tu6U+iD9UCmQvYXf3tgkWi6FLxA2cB9jFJz
0wYPqmvt0YtbiTpCAnz09ToK80VXAN9NeZJshKaUozuN6NxVAxI19W51yq161qIOROR8MRZuWBkp
Tiluk3NkZLiuh1OEXJkGgYU3EqZOiesOWXcVjgjhEOy6XgMTahk0DE9J0benrUl2Z9svogk01ZSe
qufZETJqAbHyTlq4oLUe4R71MMm0DeLtSTnOErLjGoETmWCPXTT3FsBjIUNgpCx6+DxsjX2izImY
wIxsobqcSl3guBdjn+7mR8PVdW2KAPFTdIMT2FUStbSGLLLkFoJdZ8wP4j0QSwy1CscEbTnjy5Qe
hKZM28ci02yiXrgcQyE3sQ0UPOSS2sk+QiD0gwhlzsdP5dBHpWemk2RCmMa/06EYattkRtT4/Wad
srBBwGu+OlftJJ64JmQB5Z88ztAzPRbmGFM0gDKwt6rvzFC0HVsL2Gq91/wIz+FMOc1G90mcsY4w
8ePIgaRAqaVv1NOmMaDoAi0BeGnJV2YnDsGkix30BN15gbjCEphJMn77zanPPVk9w9eq8xAmdfkp
281WLNJg/kJG920N2tYDcp249ZeaFX6iy5b1aUnZnJd8ANXpqNkqqEfogFu+w8TPjuJQIy5wYZlJ
30DFs+oYNo4rEJiOg6occkoXS65ByWxhXK8MlFDkHnktwkqSTDdV8PdsFZQKANp3CmGHul7kdZeX
/x9wwYJDYOvTpKWOw1w0nw9t5hYVAj6nH1PieGyyQvBJ8aIFcZgpJypbAV0VczN//s2wflfS0J2M
Dg0rNs5YsjXBMW7iYJW4rBn2kmT7yvsLI/5Ac5/GAbU12h5chdkB6VA918bpLyJnZ1kbhsGokWfv
PHnEPzFeFZ4HgpnOmj7Rdv69XmV4ngJ4ncogky/8qhl26OhzPLrCUXFKU3xa94793+Wlp54U3dHp
XvhMWM0n4Tze0U8rGL2eS1pGg9AvqKMLU524zww26QcsU2E2g10w2WmR5eZ4bpI2FHCMsfRm0+MK
aLuEpRSqp+6txIGfAcE1FRArybhd5W3BCVW+R9hiXvwJ2D4a1eOrRXMApzo0D6hF4CUU1Jb0cI/s
ReXC0GjablKYsv+mQuCYS3XORUEQBahU+ZcGhUmga+wilPI6uB+GZyv7B8A0F0cgq0xOrGNuN6qL
Fx21KLTMura38KQRkx3nc0sOV6FAsIowzuhw5kxQL/rPsf7ycd53sNCIycq3iv5sn5oKsyTnNe8L
UjWGQFV4ZyXRcFl5B6L3ekJnHC1fk//nahWj2C5bugeuD1YLAPFKy/uZnMDLUquq7lkpOpjoYtFt
MAwwtlTbrjf71VxDST5e+N/1J2dAx3PTNFTIxjMQUA/LllUGm8L2rO1NCkFLVtBIEP/imYxcmebl
WHX4q29T/dLxFoc9mtq73pm2X9l1gZH+8SKikQIJyraP74w3skdZov8Eu81gepNIbKz8OLzl+uuR
xKz4U2t2x6+tc9BLG8ZT4ALYX7v6M1YqtUQhYKIuXVubPJBrQhEd/5kYMNXmBVKwKKjivCn4iiiJ
kQVPIYP33DsZskvMT0ACvUHRzlS5qE03wQ2jI9S7Nd+ZL8B0cxqKWqZtw/lYAwPoHzkczI0yfWGJ
LbVSkrDWSKhFPWGC1//lNogz6MVknXk6OoZTMAYQMPOUl4Hqsvsp4Vaezyr6zYfjmhITU6GqeWoB
V0Gr4R3A4TgfOo9Ro3In03gMyoTN62osiwD06IKO0lG434FrYHZaAMVKNGO2r0f7IFABYQG2vIzr
ywBl/cwygoiN2S0Ki5i1P6Vb4naqlYfHBmD3RXWn7SKn7bpTkS8yhoZnU7G3YgT0/RAdN3nFT4sW
VZunBXctYhWvJMB+kigfrSTNCHZA8IdzGmFLOtl+ntPUEMyBYh+Y4UBnfCfqnxYOaFPghX0ORIWL
LLfnDkqDbm0h7/06lmMO3JqSNqB9COSYEPTCZyqJxFqiJx87LwEu6CfjLKDloGftf6eO4JvubjL/
pKlxxo5r9N3W81R5q9ebEc4ntOPpnuHxwjfk9mF/qQ8+jer7wuCfcLJMpOLG4bNBamcZkynZRhRR
SCkZqgeLAXd5uKqL5nM1Frew/FJy82I1+B5c0qvvlj/HfiE9NN+ViCYWZGV1U02t1OZA1ySHKIu9
tKQACGStwH79DyWWlBgTGTNOcVMrnIQsZVYnLdw64vWc2KeD20tAfsI4H++WgMeCZG2AgZwJQT6O
mO9EnDmvBJQJstSgoe+vxSRgXVGNYn+t0WTexgo9a26ySQ8W4w8t6XJX6Gh94il3nZuAIAqhuFFb
PjJQGBZUJ2Zx5NFriH6n4IxixaW/tFowrqOYfhRzHmLwliZ8QCclGvNFy36QTS4EFyPUGY7a1xUi
Y57pIJf4bguKMIGEsxUqcZ7XXyJBJnLVCPiTePyhw80P3wD6f5CIZZZxshTR8oiXBV+HFhpZqfql
sXMm4osOGcT9xGg+PvgPOy3/ElSYaPnk4XMIL1Zvn8vaSdUtkJLoopbFSh7fqPd7CVsXsjBHA0tj
fCidIUtIlSCLpeDC0wJDyqKojK0PnQmddiD0iSyQmzbqcpNncCN60jUo8CXOI+7FBVMaHunwV/tC
8FADStseZQyEc47q0iVce7d1eCVxWSVyR94AeuSk8ygUSzU6KR4EH843Q4U9mE/oWH5rGV9/pXtP
EQXZHVEiTCEpAVkfYBDLIhPgfajWtumJ4FWQuHqoCyH++i1EZkWk6P7LdW+3dBhp2PMQuCv952/r
gSpSAk0cLDMbbXey3s4QJ8NAvrFE/Q3sLHcvFC/d0Bz54dU/S2+y8o+jihRTml6aty0ZZzUsxP4c
/r423WIcH0KPtbMs0qdrFq3pcqyBtIceI5RynsjQ4ADyXtgCJuvWQYhLQEi5u8KRPX7H/SQKrQqw
eHTvFKMXZIhhe3UppDt49aY22IDx9c764eyS9+g1p/FVpznZXRgL140Nl7qbVvTEPjvB4bzmb9i1
s3+ambxf3glR0CBQK/svEDfzFdzsge/FYBuMhwzLx6btu8LMH4O5+6xKbOmLdubzPoTaTHDI7IxN
Ro/TGJaHYoZfhYBYEJw5TSivHwF2lFkZhgooac4bkZqFZWi6Dt704ZKQRImtibcUFMxaZzvTCzP5
qNENAGrlXjwwrv2/bTtYXG63FeI5E0cTBMMujy18Fd1Y9685c/vPVlD6Z9Nc+h0doDkUzchOk1I/
k3I9gg6Gsx/MsxqDr2HtaQnq3Kll4uUm1FX4C/XljgezjiGg9nVHbIk4TFAoaDcB3CCVOdWAizzh
7UpNc+mckLSzA6Hb1DCEhw6/kVLJKkKf+Jgb5zX7Oq1C963BwVzislvKf6UBLkGfi9n+tIYm1xB0
ZpiaNjs6prRm6ixU7o2hxObdhW6eVczfQvlLetn7g63cWc2DMkeksB9oBX5DUedcK8o3o8x03FZ8
/aeqA4iMDHEXjODVOdSQtDjl91RleJSPaw+DFQRdvyJMIiQR4jfPUZXqIsBJslmNS2xWPDxbNLUO
NFm/03oOnxALaOToADOTmRY5jQSrd4a4qAYbPGbe00XQTwyjg9/dUyZ5NGniQ3m1O7T4lNAH+n4v
npwHqpW9NY7Aneh0Y8UJouYRf9qgDJa0yQsC5c5/ZDdA+XaPgNgMR/xZzYZEHLIAIf4AEe/mjehP
tRJyXWDfVR3un7RFaGsdzCmsDQ97ciXjL3EtnS/t8mNOmsFiDy0eU8prYzIqPCfTXgBVruWjG44c
7rUX6PVnnm6dBX/GW0aQR8X+7+k27EPxYKtqGwEvTmNaSeC+bbMqTQj/5fmh5ULc+2AenKkjCfzm
vvqmVUYUf2bRidsYo7ubKWEkK62Lv17H777j8ErD1J/CBNw565HU11ig8MqBI775Js/BP658Wiww
vAD88MBLUgjukqbDsZfm/o03HBwsICjp3NpJYljROop8vxah22WtrfW8Q6TWt9egM7fBKhm6Thal
dGBBioEzvQy9QOchYrpDzh1b3HSbt1y1SM/Q03LXR5u38GJ/pyu8JqSH0o2X8NkEE2cGNlO5/zXT
CkrVB/YkARVkU5qBxbaJo5yhveGXIAjqsHFaEjqG1vK6D/0K1dyvxsors59hYLrOP8cr75xQtVMn
eOKHLqwNLw0gSoZmkl5ivieoPRWxqZxDNvObWibuGs8bav5um0/GIzSWq1s5hDQJKOA22EYyJj6H
WWC0zn5S6k7LyK6JaWc2GnxxZDRlfthN4f+pbvEk7SeeyapgxK4PZNeOP5dwoX5y13XNeFQ3H83P
5zrjotmB9Ld20F7ai3sOztnLedvEjEC7o4X4NrYNYFkO9Z90D9taj4N9Ca8HvytAKwOu4iyxwXNo
k3qtcVyl777wQBpIx178oVSOvSGUSYi5VseXtox6WASBbkmFaKDt03wdZRXPKT/0xaRpArZBzKX8
vydOfOkyj3oopznvBdGbqXcYVjlBpPQtJLqfO+6QQNTJWhJc8XTNUJdvoLLKaYqbcbgVxv16x50r
fl699o/s6bkpLUcNbstlyyLxjrzDU4Wz9Xc5trUy6S/dqdHJCuXM2wvJxbVonodR1juBLkufSfIj
e4j0pLrsTRRLbLpS+aqO7OS8L8rctkvS0ctosrz2RHYVcFdQRA/zfMNIlL73HKuFontc2u1QDShF
g5jq++wPLfCFNfKooQsS0u1eXaW6oc/32aXrXsaZugQM7xj92yc6abP0k2zmu0eKxYZIcJzQFhSE
0BS+xJdvBR63VRBo/hd5KB2Lglncy6uYMONxukP3az9RzUauFgCdFJA2lf9TdvQVenCF5ChexaN8
fgWzSKrq2nmzBa81TAlSFqJJVGgdN5TteCDKPTSFmeMyDAfw39zRTo7oPMWZ4N5gaUgaxqxrUWHD
fKFytYUxsSY9ynfBhF5y6gRCOaGzwGbTEw0J7TMuUD9nHmD470bX9LqN11hOS9VAsiezB8eUDSSB
iCB48NdMJdm3sqT6LKT4D0gjtMziwn4TSKbnGDAjuejn+4EgaiPSFEHzw1AUFh8kfOzPIKH29qyi
D021mbE7pgO9enL57+mkHouIRZHiIkQZHuNGM6HtmWQx+UTaGwdfVev7QqAxWeb1mjNlTzVFy2Kp
bfGgN3vomFiKtieRGFWmY+nYxF1PaFUJ8cUHtG4ydptYM8pf+O2/1GHjAbwT+D8Cy6g7C/QcPMTD
zn6f8ZU7bJpJJEPY3ZGiKYsmdP9W5Xpn3MEzACcB5r1kRhT8Xg5eaYt0/04wFrVZbVtG+bssbq5o
7+08S2bkgUP864KWtj0yN/z7evRDX9Ow/27ewQ+vc3Q6CxrqNFLWxg/D6KkX4pxBQj3jlL0na/v7
mrt96R+5lqfamj/+aIWzSBrsxb2REbFiH/ZSC/3vJ4tWnqIg8DTAM5Oz06J8oT9IdthJjKaur+Q1
Fa/i1sUsetU+aVSgpepq7vO2GJrcCA++C3+5Bduhvd0b9xc4xLUNJrBAKzWMqsceLuoSd62sjV4X
sUraeewXXpHgWCc9Z9kyHTWRKYO4M2iYOjdtFF27tAyzm28JwwRqOCvZG4qsJelEcsk0klFtSp4o
HFA5p4Zj7dcOGdg5zSc4PqS04YeHETZ0d6VWuABKdRB/pw1+xu1isMMwkYxcJE7TaW/L/ko1qaiA
1GaM/8ZrV6D6DFLFDINbb/6Enzk9Z7XA+n1hqb5Yb10Gy/TFMQhSP3mckawQ6rxWTaN1eAbgdHjB
Ugcd9gcikJ4hnWMlJDkCDapG0MpktHL39PBa5H95T//T7BGiP+EeHBIRHvbHn753wHPGT0H11nxd
uiktanL8ZAaiSuaLRoPT9hylYZk3gnQoxzTCbr8/Awe2LoDoSHKTVB2GLbSC7es3aE/X2oe71jlK
+KUpMJQ0JM42OwEf2KrOEPHeDF3XrJsfHdoxD3sEv4msQzTFEJ5MteIwuZPKXPr4PcyVUDM4rTm6
H4SrNDLQjW04SRq0KYqaaaVV4tRDFn04GCUOsl9AxROzkiHp7oCEY07rOVL7RNxXv6Tv3QsEdcUD
tBFlRv0O0lWknZRA0SJD7F3jRGcQb0yelQSApaOtVMV/YdpUamNnjHOAF/+6Mq/u+zU9IfZApaJT
OC6D5fMc93Ait2CeIzKdddgkrcONJcSQwXbg+jm3Yb/1HHFWd03krLt7hJOnF8eFQfvUUmBHomBN
jSfSUV4vttwfYfVuMkFywNo6eEJeW6X9zUl/Ab2wiRD0eBY4M3bRoAUNtRj/R4jQcozZfUrguZ2z
OO9axr9jf1Gx0imbGMFXSBfQW6P6aL1bmhI2dTlYrDXacAWnjnn2q15V1h175x4iPrVM8dG2SFJC
CbQKBJpled6XI1CAf/ouBYlUSzWYoAX+azSuh7XoaAvM3HBO7jeQzeyVv3hM2VtEPszdmdSAtxh0
249LY5eRScrjAfFu0WOtdc7mm/oNyGLKRcvsnsASBchV7ScMfCbcB/TpSule/5rPeaYxNpST2apZ
HR11sNyG9SCjOq4Ij5xQSNo3glJ+tulIEzyTbyug45GJT8DQis7LdW1aP2f9OkX2gsu9cz6XpJ8p
AhnKN4gqRbNeVfrkVxxwUphWbeaiEOyR00FmvYg0MSJCj6KOUHS0VfvNJtT80mE8WMPdqcfYyryF
RiZ+8yxa35fa7edN2WiKLdpfj1FPkElaEUk/sWdKuJSSoXu1+GjUY426v/A5VHa+xaorjWEBFSH2
ej5LeLTZUxyAHRL+XLCoBM1aB50jWVWAIMLXZnEIVqf9vW0KCzg/4FU3FCueN0aXiN2pkaOyx3QH
wgGkQh1YUb9UnuItKi8IJbxtnYrdBnJ7KtVKKbyt6RqGdmpkLhb73UnAV6sWgeBYKLDujzDv8kq1
PE8nmhHA9/P2VB3/U1dTKAE0/S2m026KkO4dWD319QV2rmJPEG9ZhX8hNPNGSDgf8SJPLsMI0ss0
jWL5hQgy+tM6DrD38uCWsj/JPjfF+aiGqfFMddSkQTKjF4fIfu03BXv+c3/JcFJMCSR8EClc7y9Q
YZUvdJ6X4Rawxu+bOjGgoHA7c1B7r9pXmfvt8ljAFb3KqFsQNrQ/3zBNWSla8rlCR6PtDH2jj8Sx
E83yL+lpl4mXflbKznjdy02ANU9h5FFtT6aouyySHm/NBBL/l8tCN/rZ4cSV5wdCVdMJk/b6ojev
P+ItvwO4/F1TgtFI1QTob92rCF/hQofBnZwWWkWi17ZTaHn6q12L08lGortdKJxH1z12Hn5jqQ04
3zEL7gnyzvTRWg3oC+bQxqq3jKsdns5fbtaZQfL8tu2d5MsBr5iXX7oilEsgGMcIyldK4WTn/ooF
ROJ17THEtPPFPQ8gUqP2qad7e7827q1M09rRlsO2pezgXJerGUAMz0c8qDFsBYXEQ2VUrAlRtsv1
d7U92yRIe9cZ0Wf5RL6YdoPpaSSUI2jsQ7FrgDt3fdula0X+nbJGMPgUNRQ89fIDzmm/GZdEAPtF
jeuqnHrO5ywICOlvZjqcpTAZRx+8lFEUjF7yKCuCuq47XablyrTWs/D/RNQJz4yJGhCm1CBW9+fD
+DaQBtKgM0lP41mIBCq6NrHU3/QB/TEXfU4PWAuYEuU+H31R9axrEJ8NnF2/vKFhb7gCI5LEDFn0
OOhrd2DwlrEk8eyfw58TiwLzyhJDZu/GWr3+F+dmxoYNGS9NzsrOy8hNgqF/8PtVagGhmx86Gr7p
SuBFXqa6br/cgJZVdoW+ugLLr27Z0c4m73cv7tFL/HdgVBOi1DQs79rAbGmWECFOQlYZOhgcJ8Ti
F3/08xhSEoLOOoBCpl0r5Z4kjBt1ATpJFaqwEMqDPJZ6o2E9FrLpXlaxQurL2o5EuFl6jfg3NIpp
x/bV86e/MUB60UgUk2fC/sHucyWmIkT4TsE4vO1qrApE722Toj19r+paQT2ouLShEw19Ny5wV0G5
o6J2fUXRpJXPAfvHucBKRtag66HMEp4hg3DAuEHX3/wU1QlIxzSfnp+xXt4jHcNB/GcwYAUdeUMj
PimfyuSqquldcpeZUWg0uOXA3tdB3+bizyH6Y58mwKFB3Rtx5dhguUokpDTmAmbhX312ybqTBW8M
zSdQAHp6v7d2/S+1bYinm1PxfvLq2aa7AEiV+6sAuBYWL5oGN3xWkP+BBIgUieWTIX1eXMumYijQ
ZWOumPUrDSsVZOO+B+3WuQCQ4bBgg8IUVhkPHIa2Hlt8P+1reOZ+CLzHPhEoRu6blnnhW/MgU9xM
+4u5ltAYlL3trPy4eBY6uhl71yu80PhP9rIN611dRWOOch/kiczwK/3uGMWuCAtnzcr+N+N4RaiC
lwM4mumaxF2nVt+JjUUGQ7bFeVGR8UsnDAOufT6H41Zq0wbEDBCgNdbGuG5O0WVos7SAvaFB3Tx1
zd400qVjwvk++7hWo8JIuyC5kpictI2LmdcfBMdyFdJF4qdcg1XtGTioEulAw7NXjCYH4IzeoyVL
Eah/42RV/QGDTFVKM3vBXkpdqPjet8FMSjC/BaYnjOG6rnKYGAsexbplj6dohJLzEi3Ni8CUyB49
xcgI+JhxNnAc+N7g6Os4GGDv3Xv0oXirc2GpqNSHNLU0jxKyUjKnpyw1FoKaRFfkG3Al7UBku28x
zcXSBNmtD9GfppCWS5j6yVy/sGpBZcrQl4TZ/1MTkK5s299c48OQCXVNcb8CgrqCkYxOJ9Enpd/+
ofyynsWIgrTrhoXrslCFxvgiwUyHn8j1+jwzKL1kPa/1lh6cF3g73bMmFpbZTVQg/aQY0S2e2AG8
8vzKGBAHCXmxbofyALz6MPDmZNAZ0WbdRJsBWM/IW6Wg5P3INpKNnmAxa+T1O5riSmfweAm6eRtK
n92xsvJn6/+2AcvSfRxi+d9Y6jsAWzSDeAcLQiJsWKojdngWRvZPx3QGj9VXLrL060Ib/Usk6AHp
C1FPQc1H4Miwj0QZmdvnJ5Av4CgDJiTHsL219QPkNTG8T/9syBFczQvUL6w/8F3+CcWoSehEiH4d
tIfeYmII6FaxXv+Msfe9s6HQ3e8L5xmVcR/MouW470mOHaEHMjPrgbFvqHLdtWd0T8v1GhibOQ6Q
dQdcwVz54w+QglJwIrDIz8vntbBRY73xd0i/PVVZcNo3cCBhu8Cneo+fCHHVM/fQadvfB3JAjjOC
5JVL/IhzX1KpaDLUz1gckOBZJPYl8h825ilewcc6n4DxITMC+6424y0XfXRJe7XyMQkg+4KSCaVm
q6mafiKAfQ2FLU14HZehw/C/RwlXWKKnte18p9sqnhxVF2kjHPPLfh8CIND/V1I3CbdJCElGa7dP
PFpdXnlvaPtsbFlDLMtO9CRk86r3nG6/bGxOCJ7gnNgt2+NjB47a+ZerwRPX1jLV0YcTQ5Nhk61o
cJl6vizulLUMJWDZRZdHE40wmkSOvRLouDcc7MASS4drGANK7UkX8kcy+yJOJUVRUO95DG3fp81V
MlyFviIXYkFEYLK2D3jMaJo5L+vsXMruGlKgZ0WZ4cQJHHczwMuLudAY5jZQwA9s5hoIgq8U3LU4
sZMhbOrDeK1a4vKKnaa3OvVvgg8rxiLkhrZcyfnvoZ9BrXlPO8ovGCWOQkI+tyHfiMHNHxOAycZo
CxnNyQflddMxrdbFBaoXp/n48E/jraEZfe8MtWDe42EO5M6VvKwIFUGFvARQDLsBZRIzr6kUf0v7
jd9wCEydGZqq7DGGYQeCK4Mqq81L6XaZ56vKwS64e1Ij1fedEdBbty9sVKEXfEzd2xNcIp1u+D2J
QzhQFITkNTIqPA8/WkiAbYaw3ZXepX8zZFPuZ9o5VTmPa1ApO8ErQUHH4Xu01D8S5aiV1JW1j08O
V9nixD2Wshe+WHzti8hzlk0tlEv0ZfJHkUmZ/4mdqWHFBe6VY63WLce/ACf9uN0/LTdw/tSEq4of
aiyfF7kgsXUOlXYODUAhxRQDx9PhjarRvwa8o9WNxzqzyq4AV2V35RM6TNnLobVqb382xsPHnzVw
SbOFtVAJVhazSIiIkriSAG6Cakgj4wQbKqOWaRk3kT6aEpi8RC9nYX9oLKeGm1JAU88+Mquj9W8R
0/VDBHMFGVRfnCvBmRDQ+BxYRhHy/6R061Pmrn0THG6MfC0NnazFgUHxchryjIWoOgdGhoPjHAQY
ImZzClZECZ0JDtjrVkoyRoTSv8rxs3Iz6egJTrVZbsNO2+Fug2QaX15cDCeA7c9qUj7J8kocUhAY
jhZroWv0YFQxIsA8BMF/oCtUgcit2a62otfyMIRu4dtHECDqCwnxnDTJ3vrpM37EvFl2BRun9+Yo
HntVLrhNhFlvBTJGXbGQsmqcBpmdCDiHzJFxk41/o6FdYC6MoBRw0OF+yPIhhv8rS42ZAcoyvxd8
vExV/qQw8FDcHUhgkfUlSweya1s7Nnp7XwXNKs6qtOLzGDq+Eejsr1CWb9A3yWPbEPVkfffLbRTq
IxEcl6Zt3y98OjL+FzBML/pVE8w1RMpcEjPddVWVfZUod1TT0VQryyxqM+C0AVeaVWhBdT0TXfcC
9gkauzfSayF9ot4Vk1pTRdogmF3cn/vP4VLnMZBH+pLOo9uSjnk5onnC9DwTN2Yb2LPGunmw2TwJ
GEuVk/ayfcDQRn4rGjm4au4GUemNyBecE2Rf/07hdtdO8bmKjNq4dC5XEWreHrQQm9rWNhQJSiCA
Nbs+vWhR3rVO3Ntx6WJDHBLsP3Y8ketVBrfI/YeonzkYmRBFQf6ccQ5k3Z6HpBmgM4JSTk5MxtDe
4e+x1HNy8Yn1BWrEk3bi140F+vwUqS5NC4yKfWPJm/axKHEkUvEB9RP5ry4JgMWYqOEVeShGZ78s
Cmcssl+QbcqVECtlDbnVW4gndjHh7Pctjy+dq80k4+cOQSHZl/e3fF+HAYa8XxrOHYBidSyFpyY2
mAiY2AucvZttkYb9TtZqGG3X8BOKXuHGw8MFUf4N4/ZKsHCg3SJ2ejkL4yr32fxMnHKm9Y+K7/ds
h7SMcg/2AU51ik7FrYZ5WtJjQ1r9peD6puG5uJ/oFZjI8E940/2fU4bsKWX0okDWrdYviEiA0DYG
+pPCrycZp1XirFHCWUVut25460ogXm6OQUkF+7eP28w2Y95FUaY02DMcmkaZo63Zkq/cFjYWt5JN
Yz6h6cy1VS9R94mZcDons2Nztrv8COd1GJi7mjAiHcuqSEGP8yvgrVbhhKGGaXxyVSFncY2R7Ibg
Z87tFdvzNUo76neKl0SKNMgynOkj/pU90GF/D3upLO9d/zWn393apfX5kot1Q/trvWAALIRabEeC
N5CgkCx92ahuNX+ZrVgTSJ+2GE0IytAmMLTPVZjQgFrzua3M/Vd/Rc5hSCOLoMrYqmI6TLR1V8EW
Hq4Rqh8rJE+Uq9nULRsGREE8okdsOaV9Q/KGl4CeIMiq3Igb/g4YakQaeYuD2zopaZ2DGpwwGNmG
XJnyXpmYz/nlaChXj6X+UqvXG2/MOT4hhsF24znQh3qFnEZU7be6AafBJy9rdkTgL3mN+NIb96wo
VwrEvdFZBKbUob4SR7KY3mZUW2JBmkR00uDKROnBJkYQlyc0H/xHEsFp+jEqMMk4KML5+DzD8t3A
HGLAeu5+BPilYvIwYQ7Ep4v6TO+vpdhPQ1kbEBJy43Ggf3VjgFAtKOyQhiLEhcFLtoS8FuE37Mux
yFnt7RFzJTVQe8v2ZLULI5BJSFS1zajgbc3HNrPWd8yTjqhARwWXr6wNv9CsY5gFeHXC899hV2Sm
pX2Wz7s+gk79pbFiF1dTPKrdwdJQfNqDC6f3yPvlyioXrG5JI6634NOUKAqu6Vy2NFYTH5RRJT0T
Iy81kpCzuNjR7vbkmt15h0JuOPXhb75u2mv1nYndh/N9MmQeSLHj10ktIlTnyzaC3cLJ9QY6d+eu
mX4jZZrNWbLD0WfrINVKKdgGR+KbvZmoh8kEEs/RxaalwS0G+IE9aD4+HMyYJ+GT+8v47XLAuKlz
aPDlcowzeB3Gkwwm8GlZrD50egzkHafBZ2jTpS6pHpDhWuhLwUG1AOrdl5kvADysRazSlEZIeTaM
Rw4TRUTUkvhzOBlmN0kzMyUDCt2fr2/BGCdsp0ploPoWq2dlNHi+Rc5x0tzGIhE9B0uvGQkcmAo1
/5GTVso9besEZFpBE7SJ7JP9dypPAX/oWO5nwonJJHcWjGxGsDLKnO0qYDclVjdko4jLL+Z7vaNb
vdH56RPDsRlueXU7Q+/I6xpC7KYQCPPtszXxW4Ng8FpW1VYM9kJwXuz/jAu+HljSPFXUAVycUkxi
CKTgiZe6hKlTYVwpZ2v2Snp0YD2qSn5oxX4Yg51DoxzpKNKmpcfDcxiah+Hpm0GuOD54o2xGsUHj
lenQWFF0G1YUiHt0ovJ+s+PK/F4OcW6sv6Bw4hmW6oF9L+n5WOVKM3I6OivsFD6lQvKE+KhpLGse
1itmMIgoWjTXpaCzIu5ru9PysLk6acG/mIRIHFp1PNnNTjLJbxLU4OFqWZYZl+3zumarzAP44yeT
F8zpZG4vUjuFD09YSGNMyz6oSo57WEmXDWN6pcpua0J2SyR/VlURd6/c9AkNnxwWMxAzcX2IQCtD
XgpnyMtBYAk6KMSk2hvfiws81Esn8pGSzRFHzyefDrmGWD8Nz0nCIGkALByFMsooCxcAYzVfkG3p
n/OnUQ/YlfW1oBFW2rgLZplH/9e03xwClIx00W/Nthj0LkxUnC8NXazRNlgIdIYIz31foL25Djln
5gEevVNce88nEc2OIu4LkGc4fMCaVO4hYW/g9hIcQ4chMSy2E3Kbi17lrVphmr9QZI02sU93DDWu
j+QrEF13HfAJYPRYjoz+MhAgddz6XGsFkE5qsIL5nrdsH9o3LqvS/ps4Eq05BBtRD+rM2/h1ma7c
J1e4RfdpTjOaWllHjzWmpSQVEWoUVB3hPX2CYZA5Osn0ZnNXJGoLErGsyeXhDGhUbiRG82pTf2By
poD86RBdG84KVogmIFrmn5bW6dFpl+kkHvA8Wdznc2E0yoHsE+4Ir4re9ifwQyLDL0RICwhq+6Dn
TQCiSNU9MYR0++cn+QxcZQ7Lb2rEkE3mt2oifPJzJwGdBqFc+sEG5DWO99AHQo/YpeXID0qhLLIv
IDZGMnB/O/sFAeXh1Wsu2PeizDuPbauWFOuTeMHxiRwnRJ+JJw6xolSjP3i2kuVssVIF9wB3MxWd
wNzGz959jvEHU8zXxjzCqF/J37TF4i17VlELTWkJyHUB3IZ2GBndCvBCveWHay/W/ktnsCjT0lvJ
lWKoEVdFlVlCmP7h47KVmvQILMugZ8XFt0TFeN9yAlxKSXzi2J3lfoEPMmp1C61mq6ifOtk+RSw9
r5MURetclVz7HgviQD/UyZ40GtBlzrAbbwMTSLFI6TSI9gfOxkGVZeQ42dAgNMumq9KD0vIeKKk5
gMxjpxgyjDIwgSuQxHzM/8iG71LpEJm6xohwoKBK5jD/Kn0r9xkat5MJxBRIPAEbX9qEzcfijyMk
Zz2io6XCwOXwgWeghvJuuZKj1YhEsWO51GeNfOlhuQZYZSZf6YCsSHWQMfTUS0KklgMBM4MRlXso
h98ZsMWYgZELRYZuxKR711hZZSRGPODWe1CobXRZNWRGfj34rFFQTUGHUz1Z/5uHTRSeuiKmZbIS
WtxRAiSZeFpC9VzT0bIHQeh4HzEpZDtmDfouJN+sVBInTRMceLTSnbjozKwM72f0ETBk45t3sgIF
bdbBHJadjQjLezujzT8c4ja4btputFEtHJ/MSOM29mZUB3J0d0vvJsA8cCndk4PHDfWSxob/aO5F
Ui0h4OrizgIHnXReJB/a84ZtHGuTbUKxx8uXLLrA5oYzilkCykeAOXx+7oUJAu4PAuOgPSiU9bup
hHwEreWn8BDIQualUx6qMb/+IlkBV8ZKvXrke8ITg+8WuU2yfxc4751NMSk3xSPIbbCWVjXdCivN
zgShgbgNa4r6LOw4a2H/SoqTKX/sj7iBY+2pU3KywxhOOZEwrKPhw0OdPrbYdHropirpzunoBhuK
zK9+4q0AYuRqwJcMkyYNCO4+ehO7sTKr+a1y1NOPHI5fjSDv5FN+GHPA5FjSeu8VIFjiNZrCFGBq
0iOYGFtKEHF2JlN9sKXdrZ8ffT1YC5977BT/kHKNNPITKCLAQ8HOrk69FEx5Wbo5Cl9ZAubN8+Mf
zXFGs9ziFs/PsMr+q7TgsYrTT7irsdi4yu87bAgmmp1eUatjQ8X0cnzelqBdanKHPEuqJLS+Vd6x
I0BdOpInwmREj5X3DkF0cduAyRI07J42MhnuR4LRBEoF+2kl5VGM9dWWMVMDy12jPakntQhlpd2Z
Y8BT7i4TVelXXkYMrLHxU+uAIC4I+RYdsFGerKKGSSM/D0NJtm/viIo4y9wHYgP457XQkMyTrfS6
CHvkNmzLiWmDk0Yn6tI17ekxeV/BtfJbr7iy9iBmuGXH3PS0MGKryXbo1p1PzB8h9FNaaL1zPCvp
xrQhlxShTxs+a6OIZqa0RZwpC/dai3PSIj1zi1X7WSuXFQezczwtznlzU1uoL6eCDuYoSG9ZgC7x
VOVPzFlQ/K+mi2KVtHlXTNRQ3oJQO79PFGRKIqVKMAjnyqmYZ8E5VZT9kyG25uZecx+LgKFl14aU
xaAndwlIFH9E9eDpmDO2PPEU+BL2HTvkposb/YDNnY9200vFaqXYLljw11YjD1AxP3xWe7Vl2JtO
8iGScb7bcI6NzaT5Y/guFdeHRJcPOMt/vb2axaGlzujCIy5r7BTCBU1Aa+BtaWWwOjvCF1+K1d2w
iFyEo3ZrsHA7eEazDPKpwrGh01le+mPpmLAxz6m/roA0heJE/0fDi5YJxW+XAQbG2U3RofWNU4S/
EpOWXB27koyqLu0Cfvu6ml2tXO7OGwkAArmhEgPGE1AGznliJ9dgXeh+btK5blygJNw+5RLxD1Be
9OfkVF6RpUyJzHXdXNHrVxobbMgKTnxEIjhm4iZCUjPq07bTXgQjAFEvc6MfMWbxXHqdJomaXolC
LOL7N/dKVxKlfCmGENAFNFWvIif0gJe2yegpg9D+WlkENSkPfazgWMb/sOmC3Yuyg00ivsDhNV13
Y+/901tlDzYg/0vsI1uU+xW7IBlOeMh+F1tQ/3T+NXUkix/ajDcxWj5MYNIy6PDVNlQWAuE1D+mj
je/5YqE2zRmOK176Yo5h63g3oGHvRbR2YJzlRuAkODbO/e4mkVdX7Gak3BhKKDJzDKV9g9nAp3Hf
bUSXRTSpKwb0TDow4vw3vNsJbzPgZ/kTV/mJXxnB6yqNtxqFj/ZMQEUBj24tV/qvaDUux7d/m8t3
M7JbgZ9vl6S0MiQCwRcUE9RSlnuty/SLm09BVxtXwPlZpslkxuAclXUjxsop+D0bOchVq5VoTy9U
DcXlvFHOctF6/21xAW+9Raj3DtLY5NMUTp5CpeNVvtF/UZnsjHnpKn85BPFlRnlXRw7AgkK2RK0k
FibDLtl+AZmcusJQnlj6YHuVssaOTijOhjse7yuaqFZOvYCrQWXdcXBvGLzLmXwMJBsfLmBLRbV/
MJQNsot/0+mnKT+q/i476B0SBTMO7zf1O82EkSBzzJ+LLRaHjV2RCEZ6mSHt/vVt+ZvGfQDW8ojR
PcpZSdBh/40hHRaFatjLD5ERa6/VjSYb7ApHuEH8DAhwKmsSyEPS+3G+NG54J6qiXpiKCHAAo1WU
d4qW/VXAas24pYJ3Q57++MPu9VukbXzqNtpE1wwnGdGHhEF/xUwrrOiU4AsbQ+HF0FE5L502C69F
mrJzLImAcUXUn5qsJhD/YiqiKKRMYQXY8v7kym4bhulXKqBX/uqybYoxp51sOJCgvdG2Zt3MyVhQ
MrxmBnDxV/4tOrt8Ax05gZWiZXYSaGq9ezmFWZ48LR3hBamRbvfS5Kq91uRZ0f+VWoC2DYcWkLXb
TOJgMKu2xI7HmroUh/CzogpZx8fsbsqnu35OO4kX8aQ07QXmiHgZvVoe9rZEGaRGyroKvg/wz2Y3
95/+7tnuvPJMOO2PjivY+twdmrDG0XICGR7BWkA26xT/DvNRhOgtllwF3B7FtVN+LDEZyLk8CnP/
/DnqYduWc1TJ8pkNpOvATgTdK4Nb4LucG8TDfUyoxpU5gDKRfqwM+xhLYVztKdZub8o3qUWrz1CC
3WuyxCFFqq01W9vC0ahCKiSvetaCt9EtjpSEE0mdpZCtNIqTVr5eY/dOOOm3iUSwEDvbMPceM/S4
qK3I3yQR/uZ3GQthSPMZ9uVtKjdjzwk3psyy1miexM87eUlB5osBUn7ipaBbl4tHuTlJsbav44EV
RwMY35hjLYXAVddBrk10dj/gPMUuLJdL/oSY2F3YAJx2tXc4P+H4GPJ/UDMZloUs8fD9teETMe0d
sLgTI2UuLMDn521zQNTfRNjVP9H0y7a6Ta6fHJ1RLy/06dAzOQcJbaLasnf+6qAmwECRsrYgQns7
/o5EnJNUr+X6CdhdJHUmUrdXhD9LWJhOo1CTuNV5VsWwJwUieV3CD9lDsjP+40Br5u8kvdd5IoQr
+3sekKwCHtwqu/uIg64g6duc52WuQ1TWpk39np9Q1BgfmIa3A1HEs79rZCsFfABgMKt1j8PqBzOS
9v9C6755s+9viKAeJlVdXEV4a/zDnbm6yryA2KdMEDAqXLeYH0IlZT1JLJGWGe37dUbk1nqx9pxU
BUw5narvvvk5evMVYHE99+mIH7//1K/9bwkHPEweteFKQynC3Rauz3l8t51+V4zSSiXKKJfeN38M
aVx84Ge8lLzfMWmhFsSzJrTnr1Nsvu5dHBzo/DsLk3PDsFyKyIRQeeqWM44JwLUHaOEwNrlatzU0
ftJsjdvjU2xwwxSa5ePCzY7FW2duWlv/p9mmZeVKisttKvlC/WAb/VQBgvcLuYmXo8cVQJoZ15PT
kpvCfxv1Pc8/a1GIGwomABp99V9L1u6Cesv1O30Avzhpnz6295Qe3gXbrjIVHHfn0ZmkQ21v0OQ7
cHJMp8/QVdrdtrjGdeYcux671x0L/iu/TLzQ6XBi+2g5pryuiCR6IBb85YfekuTlrADeWr/4A06H
VcbLu2+wI5xUqrde2DbURBgAVxUOT4FhubMXU4Apl7iMP9srDMN4qSddOpJ2zJDi0B3FX+rB+mf2
8Xu4yy81my3oopBV7+zdv89VbreSYHrqyljiU1UPv5UucI8tDAhJ3ri4/ia0LuJE2B94P/13dt8y
0fJHO+EzTkeOpVvRdBq4cLIq7+YN6MYi1MNoCfi3PasZCZvcLH3lvgCjQ95XMmEOxMktaXkt45C8
3p75A/gN6CszXHirueWAsSyB4AHU3icUj7ZS02fXcHZ39CvkAV8vNcvqYnvWgx1YIWAfLUqxWInT
gC1cRYw1Xjs370q9zmo8MWwXRjEYpHEdWFCrQGU8jAU5Gl5cBVPCh4u2DbhZx1QP9OrVuxDmJw3w
PIyO+iVA2cQuy4hX2dcakwRQmyCCTyE5l7VoEYULVpSc8QoTjua92fv6ahRgXwS7IHZ7lHREfL/h
9xRYsC46lPJkUhCZPvUO1AxMbDIR9ZrRKEr4WPO2X5bTbTULjY4Lfox/KxdqtHxOpPfWscI7KINR
J/+qcyqhw6dCzCi+IeaSVF5JAk9evQlc3RMK472fYPwVK6vI5LA0nJYhewTZo2Oe/jniIyb/Xk68
y/UoQm6MSK4RRCKe0pZ7QsB9OYBjzkbozM0FGlzuGTWJpzodgFI8AeIh9M1cidVfq0poeR2mj6P7
eCZoggNyxuMOTSUr49feSDL55m7QIwKNHZv+Ud0YpRBY5QigcIH0W7c1adlmG+xFGwAKbjClmVHB
JmjRkyN+MxZbGzJi2b5Ntcz7c6uCDdCL7us0KT396hfzD4FC4PXGyXuPSDCya3xdAAZYPrgqy8lI
QRgG41HRIm+5Zu4/3Vyj9rK3GuOhm/hxCqt/bwlmuFRoa/fBDT60P2YKxKQT7oMdnITs62xaJM/h
Tnbu9ObQ2s+vIOZzTGtzcz41fG/CdHk7BbeqKuMrqtFo0cge0CHncgGMcK03em1bnFqUDQRT1Z1O
Bwvr3ODzBj+M22PIqteyjC2+5IxKjqPYSx9Je3+mKutmgMwwtJ0polJe0cfwkLMDDlGTGqkNE04w
+xiJ6b96jpuX+p6YpiNc+VJZ2fVUJxfdWcZnbKS4UjiFR9xrcUiMzR5RMOkBV8vqloogWuunkzoZ
a82hcNTEUXP2vAxDwUDV83YheucXXdlmrCuMYjNSJfnkIywRzCudAJF+VxZ9yU6Q/kZ/JxzsPRPM
14QWhPXxoLMnA1paKcUubazU62KHb5v3dj6hnsLEHlCVoP6TSLz8YifCZVZjiuARnEa5xjYmAiiF
4ffO1BMrRKVvRLXACElj3QDgNOgMF+TxFgPUoDNyKJliJ3uSj7nJRuyY+b+sBFe4dxSPW2W9QMv6
D5BUfio4NFgiWwyTYuNff0pQgbVk3iyR95+26V3uZEVUXgfKLX9Opi9dwxz2ZbYavOYC5dJ2yqQE
jwnHudqqiYEy28Bu37T85JsTvD/f+RbAbTmiIwOIJgFP+qloimrQWXWMKIdlhEEifHhcH2ePomlv
LQKHKI4Jd7sSAqyTPNxXrxPm7opICCaUapA/qiRwEBnltFOOIJHTw0M2M+FQeS0E9PYsiKr7KOFT
ksN1dd4qlWSl82qIqMMXef/wpH4YiBzssRGWFhrz3J1CQ6bMEQAgONJQ3vORXVeFrTnyzDvoJZpZ
WgAJV5RUf2YhSwyRe6zGhqYyxRfhgi7N0JXORyo7arZaCP8A9Y39x8Y0fXKGVcwz5413t3xdQEUr
qQ15fLZQMfWJ7kLdnJBuSdfiE4PFNJrHzg5wPbH76/t3TYFcfCdhafRR2sshLF+y97CTfgpZhcjc
gd91gEFEAnxf5NeEuijQWl0w7uoC5rikfNWH/DQCv7lZKc4sxzjBE8rva11ZCIY83CMgWEO4wGd5
MaqCvFszfUzt+Wv9Z5RSjdaIl4Ufe6b/0DGF7Wgkchlr4duwG7HstnSNJM/vAv/fLGNFSyF8owPD
S8DpmYN0eQ4Zxe90gVC0Mv2y4/4a1lBdx8QMDUPq+3gdI1Tcfa5HfCFpEWqEhRfBFSCnkUvX/E0o
CykS1OnGzAT14R5RvcjR27mQGeiydHAp/paXIjx3EYt2IHqIbUO/WFnOHPbsBZbf6BzEmt5TEKhn
e+4g1DRKo6ex//5tUXA+g9uqrj0J7IJUzGk/UjE4h37ozneAtWjh73Qperpf3CluITpQfN+Y+K1F
SK5PTXDS5SYQCcS/n+H0BpF0Sb4Y7heN1JYh1jruKrQw9EEibhGAmEFTrTlR7/FDpFdePLmvpIRv
geDNuEIdtehhlcBD5PU2Jki0LA+QpL5BnpHycWO6E2SCiJmVvOekd9qwbsSb4cpTdCE5WOgkIzM/
g22mIdGQn9fAKWwLret3KNoFb3WSITLJ8AmT7eC3+Kxpcpv/l/DzLB0KAqDwqzbhjHKbXU82WV9N
23o7r6UxZYXLXD2CxPmdHjnaCG7SaLLgntvb3u+ECvpLLabnJILcaEt41VW6NyB6OwNjTQNDOaTq
ujjpRdNoolHRy5m7kznbzScH8THJ+oyzL0HhR9K4jJ1YXe95J+miTprMtBR3aRom4WtRQZT2ram9
eJnSwSN286FAmCFtxERM9piJuhweIEjrbN/uI6pSUcx9356I89stdlobytIeuTONg6DJ01MXE3tI
lgvzG8CucODx8kRq2tGNV3pXMCUrZW3oYw1RXxYBWZJMq3G4wfvY6Vn0HPs6+Td0+Zros/3jcob1
cVNdxTqoGP2hIuAtJD1DxCCOkKKHTN8P6XvMY0J1bUhhYIczw0sz44uN5ZJdHTEj/s+CH08UDx2Z
6ZTq/ehiwVKdKdrkULTrtpSkCy9uoqPX2ujsMDHQFZ4f403w6bPajS2htcLG9dnk4RNFj0zfGanV
cLz222+cJhbjAWm2flrmFugjSie9IYnK8409hakp1WAfkTK885XqQeHzCLAyZM+xPfCJQVBfXJht
gthutSr42xabm20v0mp8qVeabuc9+d8s88EZneZyJAsThn/aZf1VIX+Vt0pH5w2ucLncupC1pfQ3
ZomCfjhcHMgUqJJnrWRgprJT5SqMmmVeLatPUr6/ShMjS4/9IDvhdPRTlziTmIcklq9SYvTsTZgd
jv/ni/W4MOIAcObXRTxbZ2lNIm462qpLIRPrnsl7rKj4Wtbui+Nqj9r0mYjEwHEtb9p9RusSXHPt
AFQLd6d1y0FnGalhFESv2HEFNclLdQXK+2VUa4dU1ilTZ4F3eaXF2MNuAdLQPvjJN8j0FnrXR7bp
O4HDCCFI0vDRTu3gzkZhivM5mF86Ql2NukL3JTRmNEiQA5kwPQaaCpHhUnJv/VfXctB2zWkclPCU
c7SLymflBF3iWz4W8sIshqdj/XEFqgFHoZEHqqgCHgFhWVoFkQTNS3K9PASt9qRWJlLZ4Tt+tfaI
94HbMVGXsy/mDKKzzuZQcbp0cNOCyzj7A+GoiSk3nx4ZbezYTT9aXv8pDf/lddmM7stsVyCBJUTu
n6rG99X5M4Pwz6FWSgZUaNK3p98ce0BX4vYxx8hdCUl5AAD1BVRGK+ijpcW4G2WDBgMjRptG6rq7
5gnqHDHSPciQi+p+JV2PPTlX311EJ5SpxGW3HTddNnIwlPUeqnNzOEvalZi2hpMFeCRf821TKBZi
DbrGOoI+uZTsK1VjCfqlkSVnw9JY00RVe5AFx+QSZk9fEuMtmnKq99nkNDdBcVvryBdtS5iJsYQz
eI4JvAsRGFYchSpBn9H0ELgpGInB9DiaH74NbyzFgONQyVCxYFMAH5J1mSsAIICJlD24nlQwMIOQ
Kg6EXAshpnLCJh8I6m7hcMu3ZBwGW5drpYdmhlkR9bQS0sFaiTILQ5UPCGzJI4tyb+aGVOKF1kzu
p/eNPt4iDmP8ZIGwpEPG7VUhddZD6RklJChTsoNmxZeAvpV1V57HtxgjxAsetLhTateMsCIGKVJI
vnnKbUzzF4c6BJpoPJ5vnSIwQ9q11ceGkEWolSNKx87mDRmM4JETp1gEgYY21WpAXWemJZ+Iu1iz
uazMoZn344SZEex5rhuV9BVY3rH15RE8jxQfh/5d4C2q86Udeq7LCNzyf1XDYHGWhYgHleVvxs3m
NEREVpKgXiYuSijtFh2u++l8dPk9t1s8lwefLpf5ISRu1CBknMyJEqKL6dZ17DsqitSh4x1KskdV
jk7N1/yHAumqEUPrv1rYzXTZm1FJ0AIXsxo8j793f+SLLDwA1MZPwkCnJzHyTCeCjfWoRDd0YBD3
zFlB5bgTSugUY5jbf0B/hxFazq9sKJgI3Tu4y24y62/K8vztWjCT/FJu2MWKjBdbI3JY6vYYR84l
g68Av6NbGBNIw8yYgR8KdL4vcf2tNulBjYcSnhpY7WiCdtLBuZSwbOEJCDBJKctCBNQMUPoh1L0G
FLqj/yDimqnk3fPLJTgzLHjGxS++vaoeHEvcXCSq3+XZCE5QPhcZtTBym9oVaIlaJ5/nWIeU4xF8
0xbdSrcx5e+ohl3CyUO6K3vTlf2AzERuaUHnz5PD+ZEGxJ/WYb13oPC3wo5nHsQ7KsarAxlXOXYG
kwtHyU0CQyNGZi35sfJu2RAs2zHASYPNIc1bygH+wxULaGOFqaSfK3WvZTHCDaLZMVtxXTBZgVLg
QiRUWDdJnnJ0rPxgZ2JDiEN2vLPyXuFv15M9q6za2VCEFd+Nlnh+d7yDMFQujxuPjh2P89BCb+E2
rQLK5RLfRa+ApzxBNW52qcezc02CDaMxbvq8om/Gf27ekcf8n971mz9gxXeKVRaBoPkpc4X+gNIS
kA+d6yIFi/y8gLlEKwixyP3l7HpwdxdUQICygJe13u8hT4XYfxLX+jiOSu0B4LwQKHI3YFslfmwy
Vihqh7IzLkNtVBUeYf9zFPgPjaGTLFb+VhMmgOMoUUGZwYzjkL4YBJ7/P13neWX5HNb7zrNDflTx
z9sTxCz8S76cspsxFhvIktzMwYEksipTmW2SB2xfN1qdiIFfC7beNKXa0G6DqLd1AkU6TAB6K38u
wr6dzqSa47aJ/17OUKC5suFqNcOEYsgCAPI4CmY0nQEBj1sv6RjDQ4/Th0yenzKR1Ezehx3N5eSX
W44mXDF2bpPIJWiUbGMPUinL7rrmA2ZKkX2DoMmAq5eBPpOr99R8GOD0HZJLGvJ06OjH/ITt+xT3
x2EAuN4aV6p65O9IYE/HqM2VoapBvO6qonMN7hTCV3Nko+ipm0D6sX/u9AtEqHHMZQdGCr3q7f3q
CEyYS7ot1AfxpbsmCesIzIfp32nktl7MMbLCWoVnD9486D/ocVztUgSMv9oJzkgwAYmIHUASdbLk
0KK2DfnGOTQWYLkSIXkla1deCRA6Cy53k2feeWOYEoMij+9DTxCdblzr7c8lzCqptVWLLfp1AbCa
/wc6ixf1db5IG28iSfR72rqkzKuNVEhHtdqIkaooE5v3/zVxR2fMjMNcLCkewsmE+U9fSyPzPN/H
NOt7wHUyNAHKPYcUaW6J1gL6L86o1f3jiPrUL5HAv/Rc/xbM9XN1O+uh+NcttpkTMoUk9TKt9feT
yUJTuFkHYPLGMQDZoMhEbMOaek4apfN/zIlLYWo8hW17qanCVY9v1PZG6fl3EFdM/GUWku7rlQgI
90t4Xm6rYSAysqwXIBj45kDm9DPt2fl6jQauFmVbtOOfsWW3ZpggZKeUuhB+DRX91hHFukO32aMB
SSsuSLlqkLoEjnf9/CdNQWmzO0KNjYU8GbFLVovpOYaZBAyxKZiaFc9rMlkhJCayqiChxLRD28U9
Lv5SiG7hS2RUx6OpS4PxUjad7a27esHqMl55r/nuYQhslfisOoF3/gPxv74ZTUeLggxuFild5q6d
Recwe/Q+fmKhiD6+l7iMvjP1ife7J+75JIo5fj+M4wq1KxAH/eb8+83UsWGcSgpCE7oXUuGx2AP/
ZLQnqm4eUyOmiL1Tr0IobGkUSqvdyHYuVn3KvfrRR6mPjTO1gQp0QXhJkeLevwJPunP4nvEYBTrO
YNPDolUP9xL6J/ZONuNxsJSGFeNXuLNOIKuJirI4cVZ3ubestGtxK//hA5SxZBEf36bP+oVsdK18
gg7jeUYgsLBfsrnC6tF3n+vBt9Yec4w2p9innWK26V0sJVoDvh0n89XZdxCUpJVepjnh2T54mruD
7w1CDkTJcXE4iomSoTnT+qx94I1TAUn8Pmw1r6RJqE5e+l/u8Cc0RIvm9o15ipIfb4zdFtMxGQ9+
MrIaAwFq08/FgR2563Wh5bCp2+G4fIlG5Kmf5py2nJQR6USFs7zgOv/sLfTo8+D4q+MjDLDwY+YY
x6bEM0sROVmOVrrAmX8LLOi90fyM9S+sY/sXxCiMltB6Zb6vibER87yFK0e+nIhiQ1Yh0iTNHTvh
0R94AOCxKJB0EAnZspPegZtZvS9+HU4fivTYJVwyJhKdy39Snd6yL9MsEmcTtsZwNUcjNedMXK/f
D1S7a7URTvXsOAyRWYkDy5gNxcg7fyzNGf8Go+rIhwjl/SvCidNr46MsF9ezyr3s4Rt4cyX0A0Xp
X3LuCzcZFOXx/JBGHrK9fKcSD+mz4vk6WVwNeqpC9UtMTEblDMW/1AJVvVaYTN/TYH5YRD+uukKS
k77ZJCBZ2oeQL6pp65qIXkoZSKdGeXCvMnI9c3osfbKOMWVcHTg8s6hhsWwTIH3OUKUdtocEnGBb
Yj17yGBG5aLofmC0gIck23/mtQ0S1P/Wl1/5GqeIt6zipMBFjgvuBWqk/61wGsDFkMOPSthnBIxQ
GNvzPITZ6KaQP478TWYGJU8iwIayGkaSjQhEMtzpT7LcGG7VZyyC4ZzcQGIuDYyBOko6RK5Q5b52
VTaEcjAuBIx0Gn7XBzmzTX0u8N2lmJ22FP1DJPme4GOCsbBsnidPPWzI3eVy9qEOT6jOtiX6XPHO
kxN5He6UFj0N0ZdL3wq1YHMnPjDH2rJWpG8mIauev6I9xmLJcV0F9AIlxxOPigiOHioqISshQmfi
obhU23qbsRHVvGQfYm52XyCKrv40NgKmtKD7FfA/bMmziJcpQ7TXHvB1NP1UyNR9Pcz7rQec7ERD
hcNUgWJbmmk4JjvdZxi3AkhIhP0onBC4pxHbXMMMdEoIUP3y4IX+p7ryvopPK+jC+McTMsWtrH6p
SKjtjthcy851D5i1bHGDXzzXnN0dhSscCKkycHO/DTcPC2SLxJx8D0f/D/dEfHBqMlX27xi6hQz6
P/YEGx8T8dCfH5Sl7YPsq90pQKPnUj88Rii/U6Z6yg8yDWErZkUfHPVGgH99FQTBXUdgctpsPNig
Fg9CIhPp7UOqQNd5Rcp/SEYn/nyf5Y6/Hd8MLWQfynRVc+G7slyAUyIDOE56XVkJwL+o0Hn8HVMB
sqW4FQB77CPbPwJ33W1invyhtvYW2GY3rgngTrdZdBS1O6Uk4CNyIkr6tFxrrlU5Gonx1Mg2FQ4H
CRpYBnB+G2NfGwckswcBlosw/mco8bcjlOvRc1OQTg14njoaGZ8uY/TEGit4kDxZ/XnIzr3RthaU
XMeZXnb3FIhu/G0NeIw27+bsZLois/flVbvpqfnv5IzDGpgPk8p6BHPHNqHaeEyJ1saVwrAmbUhh
EaaoIdvdFez+LRuQCgSRZSpzNmdABUiH1xdpKlIiob2wOstKIynZD4/dtLnjMbOq+PPkAj0ZamKF
3QSDlzJiNmAIN0gSN56NmJpxmx527W6rhTnuSKSgDvLJvzXk3CVN9Nxk3ILovvnqtFhdCYaTFhdC
27Aid9mHzrqhVZjnKgIMNCLXc3GosFkyknMb/nmsX0JKkr+a+LIRtB+kbvFiycf60NBbpnb9WdTk
E42OSbkYt0vzDjuhYp9u7n7GWk4le6RcikhfgrFX2nRaZXuTz71O6gw7x+SmrZ6PYyaem5rJPbH4
5/j4q2tZXibLACQTQouRt/K2sgEpUbdQlf8wGVMe2z4b2yPpILzaDBqhB73CQqsC2MaBp8VlMtld
yIzASmWk98PUfZxAlZLvT8MnwF/FksZjBNytQ+2K+xHU2EPy4Tp4usaKcBNWd0mvnLsTgU/arA0U
Vi1V2LzfVCsLxB2r1s1x2TW1sgycu4wtAtipFLUt0ZmQEOsOf5BlU/AFUi4lUk5WdYp6YnV0i9Kr
CEm2Cve68IyfCGjVWZCshKD1FL1Qz8eRV7HsMPzn95LHC4BeTDheCFugAj6ohn196gzNJ7fcyYmK
J13xSdd4JCID9xoaN/EprLwq9fd3m2C8Fh2EFCiqg4zd8xIWfDDmVhqMHIS1HXTuGYH3/zCF8I+E
+Obghwm3vNfYcm8p9cpuxiD/fnHcyD+6ghS8bZMn9+iIo+dFKxreEmEjl3c1UW9gsSeoIxIKgx1r
ySXBTkZytOR5nmmekkXbXPqBjK38mASHhA9q3qDmPWUlshJEBe3929kopuZKXYqQZxPZpjro4PuT
k8iqt9vKZ6Fq5sbbw8gXgjoMCf9w5i4EfEOghyRMpQtVJOjQD+J40v+KSNyqWolsj+Eqbj2pS6o5
o61JfPBjDa+WsOrhx8O9NBq1HzkIyQY/BKMF41BbJo5ezLNO8D2lx1cmXOWPwZtgMi82/xVtO/W9
OL4AEgdQ0D1+R38JZJYyUUKD/R6ekY59HaonnHc/YTZ3Zd/Vw0CSOWWJLln4w+vDKl6N00Ug0HRY
don8To3lOTaWkGS0sIzU/3OZ9PjkWUZfFp97ESDS3gM663eKXAh0uhENJGdoji/nU4DNcg0/ZeFo
2LG9qgeD2cCmqH6xQOzuESFSH1gsR2eO6wJIqdkrwK+UgY0QwIC7KCMad1k97NIZAzJYdc6KGVIZ
5J9JT2qLpf5wVH9a21WeD/T1oBWDNIZgSnS7mRmyyZSZXqmi99iDsC5vtIQgBPoWq4yGwUAqw1E5
U6lQkYKUgDb5mREpacctxsVGmAEj4+oCen2dkRdx7gbtsHyIYrHnrP6b2PIzkbV4SlFQwhBu9ALL
WIDcwRP6gWElo5igAP5eyhM8UTMuy+6s6gTa/h1lBwclU6MnU8QNDSnCyiIQyur8qgXtVoKfOGSM
jZzEel99T1wG26lpr4U7Z+ZHxHg8KVCkiu82/S/m6pvFlTevYw6YyaX0KvhWb0t22T3n6oOjKkzW
5tB0bOiyr/BF6OFkepwD0nnhenJl4/K8aucFFPsA0Yob8kstvE20FlO335YUX7r3x87sGEUTPM5r
NFRV4ChNjBycZUFY/64kEd+oZOunkutfqx1Ce+KnJPmwkn8lX9DIR7L78OclJLPd29RcKAdDhZda
UCgtPQIKv0iGFbF1et7p6Pa+F2alqoj9X3ezTA6OhL4XW2T2YdxewN6En/Ydf/E4KTJe45O4WWvr
F7K0NWpc5K3hKkRgdbp4HTyBiRNsqtbM+aasMK2SNp+ilOx27QJku43BwYC6ArKuNJWuYzKXsC/W
/ikRxR3NV+Q2s14Um6Cjckr1k9X+njNrlKtRzPQrrrufq9fYeyyXfVTl+5elg4hukHIXEmjl5qbK
ga/WglnNW1/cOKCOjjbaK8Aq14odBrJZzXoefvHKpMFjYvL9WX2+RXXrctl3jqIPcw5XWp4Hto3R
dFzwfR667iPU7ToEBe2ZaS7cNGPq2TlXLDCxO24VZGgKD38vSF0jUPfdsZV7o5xng7lAnsL0NRuN
qjRr5IhvyMGtg/3JlH2gD/JjoD9+d3rW3U2XrkxxwOQiRlMcr1jMcwE99RZ1WdOtzTCywEIYZ7LR
BlHsNliSXhcBdRxuEX14/AiixtGHi9kD2yyDQJIKm4PYHFC8vwTWwLABIvbsqmjbwmjHHNK3kxF3
HuII12Z2Gd4EbMUxArztnvcgTRE65iOmvAQq7xjOgA+q5/Fd6yYglHjcpQsmO4B3vIKX9J1ucZKI
UXdZAZVcPrDf6+grenuZA5jLvqucx0nJKfztvhdmJL9l5Zdo6kiUaJOmc79zHCSn4d+cs37+AVGj
eOwA6aVZkDTkq5hNNykRiwMcrFPb4kWQ9DBu5hFgKIfUcf/2Fr57+LsAyduqqBBArwQ8eLcgBn0A
knuRJ0a3OJScR3Sus50c2Q7KzRU6Nlhx2mw+MZQc2bn94TIu3tShfqkUHZVR6uKdx1+CcgkEdPRU
NpvAnqoNapsaHO0e9pBUGZ8t5TJu+mxZhoxKdv12CiPwi3Oz03mCpXp7vJ3qjOSsJDugjFGAjH2b
57bRC63O73vJaBRbj5ZGuF+xmXf6qE9mIXW9VLYqLUzKbbBqmWL7N9IWS8Tk0Jz8z4+Hc9q9cLk7
YnBCWLZRGLMFdTNK8ggsIwkyRV0SPPrPl1sNF3Jv0W4hJ1flBDHhShKD7WBBc8U3ESDrz1w2a1dv
c5Lq3fNpdBvk0xomnlDrRQkYjNcwPXJ/BqH4Rss3hF8B9xM57JbgrbHMhMHeaTJnRa0wEmlI9PLM
PyO6JCqM7Xr5S/EcQ142rrpuuzp/MQMHyQk821Ii9y+UkAgErFllFAP+9BC327Kdic9i6V//kcFr
pSVFJ4RIJU6guy5fvh/kJOVbgvJY7/fXBlb/MkBTlfb1l9x3l4/uol3tC5qeM1g4LRV0DBQ+5jql
H/s1+BO3B5ScuAua+jcpFcd9aH0Y3thCronsSz9ZUaGYvJAWWGlrv2Q32wXKXu16oXLtWbzmskdw
MVF34p7tcg/kYgZxcSNBE8en6WzWgQPWgsYYnRrrpL0Q5eMHvUlIt5NFlQBUVtn4X1tFxl9sBbES
UzA2Fuq9VRPBvRuQb1AX8KHtqZ78NI6otFqG/x1fgl68zmW4CUMaBlupqx5TWvP4gPIW6X/20JKo
5h0rViWvXHwDSkRytjdwfztiqtRT4iOOgmKkkuFUUMKozs574XZXVkFAcQWyHoTs+plaHqTEHmmv
GmnwUX+2m2WBX020MSq7E/iWj+/6M6ix0P4/oYQzUX0OiY0h6jOJgLeBbiuHF1TzKDQX7LGKlk5P
gYjByOlrq2e5dxmOacca0aWjVmCox18bz/dcwwHdTyUnlYfvjVFdQpMiBTZWq6JdHgtFjsvxc/aI
iDYizLmLjxPnXEsiVOLOM3oKZv+ihTMtK91SBAuUAKfabwYrLoIA+yyYlCv1j//WguYe/RMNlJX2
NK9WnENZwpXRg9c4ifdZmcDeqeeFTOlm4NusLv80Vq1UmPC2xtOPp+zoxYlzv4Vv/YYrTlfKyJTl
YXo60GJYYo2775ALRCVLZ+TWIhvv51CPEqHHbXZ+0fffhO2YCAIpANK55vyh6dN5o06tVVYS34Dn
GjrkKaUgk1yoQHnm18zXwVO+3J354+NqAv48ggt0AttbpfYpezlmLvniBKfpyU3qHZb25ohczDpZ
oUdX8TZNET2v65o+mddJIKG9XcsmAp/2SNqTGB6k89OssR+Ip2jGbaoRMckeCs9ZK8BFBazQllUg
kmxJl9viN84APgephLJhSRPEvVJvA5U1V4QgmzxXPqZpOadAtOFp3gzH+zYnvDo0rSfcT2OyEv9E
4CDLBjPzcwKXXrJhCc3zh1Z8GgHbP4NpgBqFhI5NDpWxkfhCoEAahfQATxsKFk8ZAQoZYsl0L4Bv
QbgdJ3Xs4CSgVPE+CAhGrsrRoB/U2bMQSCQ5HRyi/QQ/15M4mpoqZqv2uDckgBjtT/9DmDxFU0HY
JZeC961GHZselsCb5t/AHiTwLkGvLOiZ45BzMkB6W1gp3QTV6KhL5haCN2dRR5lAKhTCrSEkjRw7
TCgytPraGVSyDTat8Czco7eZIu05u64EkZUuI3K+VoSWnMLgN27vfcTGAX0s27+jPqV4PXOyrTpL
Ir0Gr6NbBlJDzyt1gB1BleV74fwcjDixWa4YmxK2ILqgbAZFMXOXEQuUAK2AmMi9uFCcQjUEHgHv
dVRzewE6YrUZ3irD3sSOHDuXWmgUiCxDGu5UELcV/nBxfjmj9ORQNAWlZ0LSN5w3xT9jSNFbVZ7O
Ps0T9DPnGjvQa8KOMzxTtD8kh23OoB5uApdNhzVlKo2D6mmw0uYxlrGJi+iZL7siqYcoh25Fldyc
M63yKsjwcUq3a0BGNCmbuMnepb1UOseQvasxhj7KGRq0XsNk6sI4c3sz6nta+/Zci3hXpz5FuTX9
L8WVwGpDCzi0iwt6+VigVc4WPdgZv9VBwZwHQkPFVJ9fEVgStdL/EhapE9tKkrR1bUfkNm9W195C
q31L52A+6AnjA+VfVJPJXVpMk5++1VfIOdhvG0Y37L9YUKYPfyettTi+q78xvFEzmVjQClOfVpKa
cjDXKYhznNEw/13UFRtV1lz8C5jos2RfeqIAEmLn7qkSjFWFFD39tvgsnymp9atCFVEWNqO00Xuu
Rday+Yu+jRNqbURpDjlwfaKKdL0Y8ygX54MoyrhHOnfTTjaYysPsVkHghACbHWhRfdwEp4JPEXBq
jBYsmcDAHdbxI70IO26IIFefsM0HqaqK8I0rNpY7JVXWikZZIH67MwjbVlzo5IZ7SZ9HwUvjjQIa
PR92igsUWqhIbiiwk7V0mUjD18cepVWW+vUKKADyOWQG7bGWdaQnf4WaUwHAN5oFt7hK3iZdZ3bd
1uQljEYNB2QaTGzAXIigm3ngAyG4qG4FUld9Zi/7wBviCMEoLRZocS1RaCOBUr9lkKjMvCDOLrnQ
FK/iIIqwHWBsQoBcfs0LF5dVrSG1YCsc0fpYHehW33U9QRFUq4LTfO52d6q5V3t9ZSgu1bK/4Bup
z4KTLh/juoG3mfPyfQrh0QrrV/fSqIQ3zGO19YS7FEIaqDiItMyOWcvtQbTDJOvcZqwgeWcvSbUj
BZXKwPK26fKpxFJ6V/sAo/k1zNKTYFVHLCc8fqsg7nVrbk83xTHbtNneFiNJ4e5wRD0cNBuzB7go
kcQx+UjsvbvTtcxL2RMbIXEDd2GrmzFPDLVfaW5FRebv1NIljzE7RRMEwe6KJ6cW2Yx9Gm1lzyGY
bvl0TpnO73y3e91qJdbYWi8wHSXZ0O4DcgyjCnWWfrBnYZEojS7XVJIYeCynH5hIdIwV+QC5OKJ3
O1M01Dw41HHPdvAMli6QV4PQ5sOBwCUKOvKb6mXgpMEtkHJ/+tOgAClKTRicK3bsvQHDr2DQca18
3WtuyalEsYJX/3KPpDBF/jRrGLRE9dXv+tTuWv4L08ZRlT1uMBtg/bniG0vSOnNUbh0NwYcSagbB
mvLEvGK5NT1qNNFJu0E8UrHaUSLqu2LJpogJ1H1WmEZOvYk5bp4QCfxfkprY6ZJx+oCiEsnQx9Qj
Ga/xTV7oEhwGDSKVKmtXHqapc99yAZxSoq/+KgTPONpyOSFv4a+xaqK8274AoWBOEYjPpuk+pUit
BDkgc8E1w2VqnCUiceQnLBO/252CDXWIBtCLpkXBVUH/XJMkIyEgZwGDXf/76m1rwzwEe+iue4Ko
JTcqY3K4Td37auhsAVMhjFHo+YcD8jbjNdCcGcjOLzL/F09LnPYgcir7NneXbg2H7CsKtfvbBW5H
r5S7pB33pXjwC0/UuMBLsmgQyPm5vSa3cLyAEtgEtZhe37udAewn2p9SlIxOUpW6HsWHZBIL1Ljj
8gkmdJGy1c2jvqINrzm+2bt+3Xo3cXk2pbWOAoBqN1I2BBcjt6NZ6WtXbuhUw6N6QeNpR7lgr9GZ
/zZeXNfuR38eeY+QQNTqOM25jn/lGVJ+jXIAy+247t+uttxxKum+PSJUTeSyJP1zMAajftwF4TyL
R8Q6w9ETWqi5b50M9veOE5PrNtEIzhvTj31H1XqoVVKa/gFg4soPwDZGCwFjpxr4Pd9UhHn1aZ++
g9SmYLgUJk4gdUKW58qpFsxHDnWhKO9M7AnUC9HSMNJdVa/15vyWoPuhf6LojEJLCnIqVmboJNjA
TqN7wXAHdeVTROzf/5zsPxsTJ94W1SMoLIzXmRhGmGfZpkplOonwXYdr2nruY+bQZQ7LJ0gC5qZX
g9Fi99wPOC6ZXeOIZAsBmY5smpKCa2H0DxslSW45UpzmJ9P/zjJYyO1MN1iivzSBSbc1yq/j6wP1
2tHJ3mOZOkVKq5WzKD/MvthdqoxBKQh+4PRHbNwFINu7Dq1wTdPz0PDiA775do0FTaK2pj/49Z4Z
bfmpK6dK9Xz/Gw9lJNfHJbTQMwSZaAosYF9UwN/xbY4a3hOa6hnzaz8b1+N23MVDHX/laP+VFV3A
t8bHtgQdlbc2Q88hj7g5oQtyofVNergJgRoqcEIH9U7C3eQU4Wmbok7QTZMikpzYsOJmevGoIrgz
YKXAof15W2DxDQyKVddZofvUGajjG9e3sfMPY8UKAkADWtcEsKs65l/ORfXU8SddD1EMo+9Rqnwf
mvjhlHS5GNFomIBg1istATFmbHWcHC+tlk5jwmVyC/wFKr1VbcDMm1DNz1Ug3fB7Id/XQrSuMQaT
XBnTrMvb7Dyr2z7zn2f6YCljbbMnhZ2Pkx6RVmKu3Rku8X9peujLcXn3QnCmOIDno2PaHw+yiOKF
HlUd/PNMr72h7EHMGL9V3vNByTJAYvOiut/bRFbTF9gYMlc4LilWppHvObtEdSjJazr5KdIM89sE
12TDhJEBjUsdBkFmKWVHAmD/1Nd+CRm2sD2FhyMhbWvK4bgiMiM36QQtAs1WPjP9ZXgW8zwlwzP1
keEhh5TBiSbhNV4RNrO9xCz6rOJFSqe5rHPa8kAej2U6xby/DQHUQ8cASceXVhi0Bv43C/t3+jmE
NUXLQH9JoF2ZTSzCBReWJXjf+/OgD5USEjXSoPu+SeukPAk03LFIKcgHhViGd13jGdex1crJPacS
z9BiHLec+0iA390coUZBJGn7W+94xGY5L9z88aNF+ccgps8ZKiicVUvf31bPxQ/5J4R5sB6Bz5Ye
MPJRrsvpoVQyoo38+SvMQK2jYBNR1NnIHn4rJoCHOtvd7kjAxvjiiTi9nNFczLCu+pd24JqLGNna
OyiClFoUhH/huCClmNlZsKZiuGJv7TFhkLKJOjr1FsYFCLBAbxY8+i2vezyzdO5oBz3bic8O4vKp
EfTo07NF2ltcR6Em7CxFRBF46nCUP6oSl8ZhOK5xkl6xYJaP3cTc1quNFY/DqZleIiiCpoqKCmem
RJ5FpWoL+4YsgscdnG7npHXM3yj5IWdoooWqFphF+dWIMH7hKattLWF8OfGCt2BotlVBKjA/VOtm
me4dlF9r59+ZEB5aMyvD+C8mJAcEwRE7qYIE5CXQys7tcaCx683po3H91oGqV8AV2pcj0RMz0tB8
kkGFSQUFJ0e1L9TIqADWyezZ/zupXaN9w9avSNfujO61BuaUUD9y8NY/M1fCtQyXrCCsWLUtyXuy
3VZ0G8zU4n59MrDJciH4Br2NxxLZx9+fuEXkdm+8SDYhxUP66XSsxgub6541wlL0rg7E/Fei1/d2
6ehTMv1u1HBy6EHpLcY7wLWM8BICL3qInUF1YMrlGPqpZsr3MYJIBkqDKRxkdSd6UEaqdN0BnQ53
dYlg4XnnTCue2CEPGBOQAycWwQNOze/2B9WTyuQ7lLn2B/rzgD3SpmT4O3xzfArbl60nyL0vbpL+
CgeTJHVwz39u8IQTOlTQlk0TJx+EzJuedxsIWBoFMRlg/fcxv5M+GW5+RtvIWlnl7uNsyzj8S6lm
63Xg/JaRmq8BSDyh96T1EnX1lu+P/Vf66fr0I4+9PR3Az8jZKHJzKOHK5NeRqj15oHMGkSdshxDl
1IV35F/ofuOMEQ6NrZMFluStwUfY6ayawGqqn0hiHD2Mb0sMfzG5eXHV92Inp6MF3uhxttMmsDBz
0/O3x8fhl3UTO0NQ6cd2xn7sbp0s9MSITUAE9MSDlkA4ddVLz/aNC4z4tNi4+2bxYIf/Jw+PN+r7
onk2tFBug1JJMUdI6GeCCE82LLL9S4YeYyHQl8Bl1R6xj3AV4A3t8jk6mKSMp9qRMBqJ+WQFpUNs
nCZ+5BJeDqoDMg66Oe/r0JDFByiPagWpwu8ZB2GmM1QOg3UGovzAZiujx24JAUFUvJo2O7ZifNop
9l3cPIpzr7LzsPVDgY2rKsxYIKPAeJSdowo5su3xTvp07rs3IY6MGJb7V+iC2mQGZE2QiBeMdboF
SRbwJV1OLW2zR9LZQCBdy8h0Or6OEjA/zM+NJ5e//NPdJTa1ed2FmeRbLlMvY0GlPhnzcf3DK+mg
VhpHHvpM7hFD83pV25qz5DhOqTUoZVdVa+33WhMGg4+Y9AdOGWpxTvTXBTzMncEY7KnoN+Ac2JVU
+ggyZdlHpFmRMDoL+/NeRKJzbOa/PyWoxrCPK16c+CbRedGwneX8Ql9Vmv74XsOOpQZiZMOoAnF/
yRTMo2L1Zf3pGurxvFgwJCEdYc78hLmc/qdRZ/HGN/eFa/1UK476Fzs3hZnJJqlQFoNVHhFUHxZC
gGvrVyGKO9Pd8shg0EGrsKahSXd+ha5dVDkH8NqbsAxevDLPmRdrhypRhWtalTe29p/UPqhs1Yag
M+ytXdrbhkw+vYFlkmo37PmgftrJ2o4fGLHNklzHIfBa2JiATx5DXS1iHsf5djCD2SeM6bABtqFz
133vHlL+IuK1CysbS9pJ24v33Iq4liEFqMCxs8hf/e+gavAVki87Xkd+/vyzckJEGJ/QhJjw0FI9
eecLrZ7FCNMp5UDBlLnAobo0BZAQK5TOYsUDzA0AvSV17TtlThybfqNyh1JikCUkbHGjBdTEmyWN
1EP5iXMTeuNNuMJaA3TZlDiAMP/E621OgDd7PKNk0e/DDC6wUWMv0O1IT8vPSUDSpSgYDwViLaYJ
LSWzLzZb3IRJQgFwryrY21uVosxBWfxs+2rtZ0W7+pCECLCtG8dIFAeuWpXN4AHsSv7lfEe0j98o
fWloQC09FWKBS/abZ4gBnHaAK/+/6i8lYCA1pqruh7oEC+ebxTKF2V94McCu2stPPntY3yV6tGuw
HNw63P6ZcDx/5nGKx8ZjqtkRHDHKKOwzuwpAHaKcTmX74kwf3XyRuB57WBq6RliRYHhMthh6aEHW
LZ+gFcnVyHIzqbvRZ0Pfsr0mRwQ8QjNYRqI39xz4VJ64juv/5MhH/GPDZtwJpaBByQYh7DIXbfmp
+DCxyuV6vL5dwtNWu8Dlsb+EupYl3dM46GUxtifE4zWJVckKh2ZRMlEsqlKYVo1ivvlZw2eluA6x
GWvkaCvP0rGiD2HkIcRKRU0fc9wS4HNvKMbd3giMJnmU+CWdFMOwUgTqmccfnxwwuzRByhSolMxj
lvyGQhhODc04wp2jbmZA6odvVLi5CE+7pjtTPf+Nt5d+oZf5w2Bqobf0Uk/7lJSqu8KCMgSDjAvY
urexUstflAM6vqes5Qk2Csv5IAg4RZuNZf5Hpm6BRRuFObaz4SP4m9LjaBn68lzRdUlI2bOLl7qo
rPL3xyfMwL+b54gnWstck8Z9QqHS4ayLT2t/xLVFSIJcwf9IKtvLn1npc2xyxFc60FGL6MikEcG7
HSeAnPvTPaS6OnTha6X0+fdNjarAOj5UlwHFL7dOTEATPH8c9Ol7r1TL2xNOShQ3TZdvqYNAQ02f
5NiqC1cr4CwkNq2kldT4okYp6iPib4mGaSuMZ+NGM/1RL0KVvuFJRNfu6z8tBPqx0PdOZL1eh6fe
em0Effs/FTF0PYOA4ZNGCA/8yWKo/FAS2H9CN6JOlH0ii7qotLwSs/Qq4o6veVC7C1l1+DpRCi9j
JPCOTIMnmMbjXCgrQAlcKu5dY8S83H6pkskuWRS162jGgxbbgQ8yr3lARK/IeW0cnjt4eubyi2V0
J28CRYwXB22BWsONHWCR8azPu/sNVqGTyvIXb1Bq+VY96N2dYzd3KDEaFuqBFSnfmL5NHCp3hLTI
h3BI2cbH4+mhqxhso4D3akzJpMYgPTpjs+QaCG3uFTI7WawbG8GhWcFjLwcarDBUl6D2n2mlBRwP
2pJ/Y7z+L30g7/R/GAimHzfy6kNk03ZUBSrM5rVlACSgqcXpfcG9LmqgGog3wphmgB4uxLULjdG8
5NS5at3OAI2FtvLV1/NZ6K7IqlEWhszUf4eomKVuz6sGm8jG3ee3HYcr1BlMeTWB0JsBpXYXRcGv
W8PaeAS78f0AcSacrkY0UY9lnvldnLqNDOiPpXloEhkeGkpLhL2SfnLO6GachXgu8nD7M1pUKpdU
IbjJiQbYFbLw6vaj2X5bNmuVhuTwH974PsJNseorMwTkV7Y7TY9R/wPc5qygaXNFj7L6Dk1JCPyr
dpLIaqxJTF6SOyFyzhJ90BwHx7fQq/kPhpA7fZ8L1MSVwDVrLCL40mdm5mKTvbyzWgd9KPX6Nyry
dw5Np0yZBtquQg2MktFhC+Ja/x0LVf7iiCKSeq+GvNstX4LVzOocvcada9OnxxaHysDfUaWyDYpD
DGAJsWfSse7JQ0138pQygSBgEb1VsIWkdrsdKy0lP6CEPt5FpDieQ6Y64OxM4KEAnpogTHdFv5Vp
KynVsuBvxBqezmIkWIiLSfzuuF0LNk/jx+spjQqpV642q1UqW2gX2zF0IDa3vAH0cpa/K1oCuuXG
PDCGXH/jc9IWpj42/1Gvqr4iQa/56uXTgLQxD/q16dP3nIlE9u33RpOnUaFrf5Ulrv+qteA/3PkT
QskyiTsybLkYqNt6qKd1e1WekccE6ynoYETkKXnliV5NnE1f9UuysZUQKkNHy1GvyPLex/ukL0z6
YJq+JDNBYBJjweBY9v0w7GtTiW30WuW15LX9KLHFXABloMSHGJS72NDcsEUPqfteDIEqxSDGpT/6
b8iti9V1COx0yRuehfn6mMIlFHPiAt519Cdp1wg43JTIL84vgVL4dg76s5I7zNRLAfaFNQuZlF37
kfF+K8Ge9RMnIyuX2RlHMyb4qNlY78ZufMHbZCzR68eYolkAK8mxRjJpdlPdVa4YRJ2hatVLuWBD
lSsp3qYOHK7dqgT9ZWjtnOhE6dXV4wYoF5ZhgEQO3htum/5PoqPMgfPY2L7zK3PE2vwKTHyPiVXZ
XWePN7F0dkrAd8SJE8qwk4kJLBsQD8VsTzTUVAfA4iLPa4ndnMnUM1XCy0Qylx9B+QiSlWO1QFqW
F9Cv757wZwZv/urvIwNEmqWfQsn1w4RKzZEksP6b2P+bJMTymKwVefMd8FEOrlDpK4lmDDfPuYqG
YjeHDzUlmYxGge8I4jOaDB0hK/MUsfuGMGzfqYlkxQxEo5JvUXlfOp8oDcpZM5EBRQyC02jN+CrJ
EvMB3Jlr6Vpm027ZJitj6fi+aAW74EXu8WJs+Nxx5rbxRqYp8/vDBC0084iltzsGwK7u5Mm110pv
2Ab9REaMPVTeSi6PTt72b/GlyZAzdmEAvKksZTgT0EqlolzWuTWdx8tAEwQDTuFFiwKXiBDgnbDQ
esyY05sJNkh8Gnb5t0HUwHkjdP3ZLiUSxnjOiUgvLNp05x9O7ZAPN7btIoprtcLCiN5r6gsA+gRa
OVOHLHiCPl4X6N+HhZUP+f0k60jF2beLwbWezpmf3sOxCiO5hUgvaMAGW33oted/aag0JKoJp5Rs
Wpe7PHK9muE9CDBMTKnLI8aQukMz+UMepVXsyellsxRhl1GssXNkOYOytQK3BNbhKP6g+JRaEhoM
TAh2RaQfeXA1Wx0Gj/8hLplsYoGZCwvK+Yd7d9nFyQDHJItEcmKPl6/9nsq0k6wuygWgtBXbwGWP
DYQ0Xjrz4+tOtTI2A6HxFt071BOyNkBR4m8JHkrr9jSaOIo1y/8YHWSBwfOtRZNAjok6vORrIGH4
MuEJAwgxaJiLJjKUpRr8MCEdE4QhwuSRGGIGWjPhryIzTyAzsWywi+YvUH+iEfYDIfcOv+ivTZvK
lk7lNytXqWmuA1uqXzHHLJ4DAjwFUWhEsq+de4uj5eXGEJgZbUxY5HQSxAN5wxdEaq1yMZybrIos
XNZtq47qBOmkHixNwdfhRvUZZgTZRcOwaNCssFWqhy3lXxCEoM9RgFxDOBTF/LUZKE5EiQk+xuUw
P4mourAtbpFoA0xRYULHlSS3h7VORdWf+gYmcFJ5J3Ata6WVqcDwBmyp9j1rVKyjr5VGk+jj5Ub+
doCCskeYtBP7ByPrFOg9a3CBrJi/1UNaB+svNrkR8pHQ/8toN+JBvfPaxlQ1fDYMWh43lBGNVvyi
Vxz6zNUq1G9oGfOdic6qNScYbQsaW/BOQ9xk7u41M2TbNwmZJCUkhTB/DlMpL4Cdwyg+aEmHclco
QNPv7iznD6BWG3pz9LusFZh0IblXl1jN0sQIb7/xxW0ofZXuTFBmubSiRIngLwHG5HJO9BeBnjpf
SDBE9cNK4HBbJtSJB1D+uL6VyQSz2pxaV46JV5pBZXLdNjK288WH6IQuLRsJVirLf70TKgxUe1cN
kBpxqmPJKaH67dRs0tqAi6uOk5fgfNcXf8wvndcPDr+90W9+da4rjD+36TkX8P9kX7K2yIQ7RD4d
5cV4V/4nYLwenAk6EJOn555XohtoA7pxRAXxnJXhWKhXIDtrmkSSaLU/c2Qc6fDbYp0PoyDwBuRK
Cnhz6XYrLN2oyZZSnbAk9uZEkSt+MC6b9zZZCYygs0AR8Nej+07D3MTHIZksk1gikxjgxqB9Egfy
81ndbxAqUeL3x3oOZrzKIvwB3tWBlii1Ab8qZDPD8WDUSz7p5dIu1nxVPnvQ15YDZCu9gaVVG7JY
/YPgdGzf0A5ZfvmFSvTf3tajs4bYDxmyNZVnbnqEeYvvtFF4wW1Uxrpt5fV0nbQXNbhPZK+EwaHv
Ukw27/bmxpOqyCJtOjCBITqFziflZSq9mBoS2uDwQVT97Uk5E/d8Cw2az09BYuwez4ytZi9uPT/f
fayLbXiT5R1hVVN8yjMsYMvuIJXFvLs2eai6uuvcdCdtWp4kwvhN99CQRCHsSzPmx7zvTc4paIbp
zFKaMAnM6axNCtQjvK7aqQJcpdKW8426WSo1AH6rwdDU1eCiO4lIZ/szT0u3WEe7k1JjKg8pInX3
+h3r0pD8rJUKZGQfQnOo10W2kiK/KZ+4TWPCAPwnwhDII7zKQVXP43YXBmz33I68nYFQ4IqTJdqx
cu7ynBRJkSvtxuM5tHiWv/2yiCkG5+HSzSZJufjIF7Q/owtcT+Wzifv9lErBpEncw0ZFye5qwFp0
8s6Wvw9ULxQ2FqK22SBkr1eRVTr8CVJ79ShNpi2Stvz3TFRMd0S4Uox8vB5d8nLt5iMQA9tQ3DOB
kXdoHgGmoDYfi54P3g5ZbwQYQQPSu9LMnUqNf8J8BTagIXxgdM/7M8mQXN/O/qQ3JhTT8cUGO7Q9
i+uV+UM6D1CfClQJ1/CpSvXNfbN4DrxJGKB0Zo/U2uM9zDyzYRs0paj9VOyNOH0xwbMJACKpjXEA
I+tdoKL/H6wHfcTElVV81sdsfjM5yv2Uq7muqmREHSavNxjh3PqV5G8UiXMpgPfmgufwGS47N7aV
kjUv9GnKxdnie6L4Ck17TdrEqCKjOr3fDIlpHzZ8sdsAHd77Ejjqlbk4sbQd7DbzWBYQ3SXRupQo
18/3mgehoqp90lQveiiuW8m89PABChoOsy+tgQawsVjBN1nGz74INukBc9x9OiC44eJEmj28eAhT
BVbS9ERKIwtCsGHls0N/76pqNCZ3ikDDCYuXXENO5+pt+QKtK2dnEapMpFg7ZrUVfCRX/LqWhHvr
gznw3IiPfXmh2+aFvEM0nIaoZb2L0z9z+eARIHfX4WXYtMctEqQUIPVpIxQRvOq/dmB+a3yUI4sk
/zSTNe9DgGEOCkWLQUf0ClIgn9tqYVlpBEZhiyEiOM3ACCNYz4zvGBSpAcGUTus81hGVCLoDwhTl
cRbcWwMDGIFAgzGvrWg0B0PXG6FVdSUzs/O0W7+R2ICG5GPNb8HpvsnUtDQA25lxvIqW6d6uU+j3
/GLnpITMDYDvRq5TG5UfxcbMI6hp/Eb7Yd185SXq60JPykjBDrVfUX37+3VLYM/F8tAXsZrfvFyQ
Ox9dz0NN0Srn6f/J5jvOi6LpsqlVw74sXdEgBK4/X6Pi3jMDXG/SLYyNz2GyF79Jkvf3sxJ8n/Tr
Y4uwlIPMoo5qruFAa64KyYylN80hgutbNZ/PLwdcOoyxuIfF+mDAt9aa88OD2zGCQQ2V6EcxgLx4
pd1ypIpQvnFDenoD6d7aAleiafsmnny+EyQ4w6bsbiyncMQbYlW9HXuq0IOWLIaelLiXwrvad7cq
4JqV1hA3a73mZbNgcn10OrMok3Y0jpcag9l6+OJhvWtm7G2gYZUJblHDegywKkX4j/9OObS0SPLo
DG94JJZ3xGcLC9+qQ+mLninR3P7DpTAJFd7DcaZK6PyY1ejT9RCp531uquoKyb3gEzDL8xVOIFZg
ZHgOnUvjesJZwJZ0fvq9Zg6xT1hs0eAo+u5w/F0fU64Xuth3lHb/mKO0qAjwX/mPtImonI5KwgqR
wU+3azbK/AxULp81b4Xq+HDhSbR+h+jQLtNlk0k2SkPJcYNp8x8F1/1fyxOMKIUNxJLEWxZKmUwA
hoclhJvfwMnL/Rr0Uvh9YbQ7aJ8s2VeLNq31ojPk3plhzKIhr49xlf/CtboUXsLvCdrySw4P5XXh
kUJGss/vqQcex9Hk/4Ny6Ey8+oaGMzZpnz3LKZLSsHkWE2l5mD8f1R6HhypKZQ7CT+FP1tvKVXSZ
OkpEXWMrhT+TJEfidU1d/DCdGQu70PI/BVhOJmPWjJZJW0lKwl72FyD7qL2nyVT+i9qjpwgOYQMq
grJkRBKMEVK+y0ZWqLC/Sf4FdMvmyEHIAExyS673DdPbV5SH9uLtJiyijH/54MGllOxkUNdfdits
X+akapMqp+qha8/OAsBzSDWdp1qrXjJsss2H60mjhxkkoFQwX1NjLAr5ueSbx8O3QdEoqAINSKTf
lACBR29JiRWrLqjfCU+b/vQcbRQhQJK4/iZkzoAS6eQGSefOAE4k6EtRWrDHU8T2/XR8oY/eWcJ0
jl9T1CsQVDmd400qzNl/vbFepy48epCRlkWcRc0uel8vxhtaDoyz6dhoZoMU35xY3F5Z8cbRo8rG
EhGyl6HgwWWHsvFMwAaIXJ8hFqKr77Kgo6vNZPxKmiYcZYTBic3VJiphy9gyLC0c/eOnnZRiiplJ
eaRDRE3mdb/VYbBz/Q2X7c7jM+KytLwn68eZXKfYjj0Ua97DKufESPZ02uqW4INH3VOOTy8FsSzB
NK2+M2+HZRnE4y7xduNxwdz76eyunS9+EJ4ptGEoQtYeVrkePK8HGTqNvlruGQA/iBX31EwDN1Rr
54Mr9m7ClZTUYJiCPD+XzuuhvacRb0fJqMDMVYxDv8nKsZ5XFJaBKsHq5G3SVuV8qWn3+PKjGwMN
pDVdtFHbZurZLnT3vwNK8EamxRWjgzK2ZvPjlDbMX0DvLF+1bL/r5eMIdZPEBRZLkZfljnP6ij8K
mqswKPr82OwgCX0tco2aN84TUsvO+lYKUjkAHZkL/ZLOBCsrz/1aFar9AJ5J05LIvW8eeFXGzB9q
UTJ8GUfW/LELmaQQKEhRSK/9neBDZr8SJdF7QY8E3CMjQ3NtlWPNaWixE+nWOZN37U5e0strlmWg
gHmnslwepU5+PwKMSA6487UZgZIdiOxIqmA7bGFBRuwU9NpukUBwgtz8GOQd+jk5LfbCCM2tB/ry
r1xQxNBBQpWc99pa9XMlo0OaCzgrE1MsvbtV+08saZ15n9r78pIa6POizEi5Sk0Kv9Kt6MfEycA+
AnbwPckwH6agwlei+rG72PrKm4UGIYeNeGH7xlAS6Jf/hVqkR2cosbTqTGLf7F05uti+TXkQKkLN
u+wG4v+4Rwey/4rG6NYNBapItC13ZFBYtoJgpy67URJDnZ/hBnK5oyigs+gLRzgmLW/QU909Vj6h
DQqiQq20m5Odb/aw2rUdCouUzoNsRs2rhh2E62zn2oChNRUpq3ZGEJXaHxHccyjQ7BOFqNmhTsZY
8jJOn1HfVi7YcVzgoOtMcsys8ASCjaCYgnegmRbLCiXo9pNDCODbAJvnc97SijKSk0QhDJHz47DK
uaKZsd6rpiX5u0JjwPnKB9iczYxHJ9PToOhpbSvP8qeDK5yekHPKdIeAz2Cq29dVE3cH7URSDZPf
i11yAZSVqg4bG5qShda3bFlir4jv5EA0KnEpW84RYbektAGpJKnt/Y+MumUls0Z+tO8M+TrnN+Fd
kmdR9NWj8Y7IhJFTZdkXf0otH+JG8Ny+YamfGKok5iwzgDPqLA3rN98kdj06ivM4foNIJmDlcSM1
ruXGJM8h6ebNAdcT5gpT10i4suWQE1IQ9+kMf0nLsv4veocubTLXWwYps1aODZC3aAlMMCL9vCS4
cIead+qRzkBYMQxtAtch20n2nzaFYD27OhPCs/WyJZIBuluVpUll/oH5AT3FoHlsOoFQ2k4qwPBZ
0oh6e4oERqR6LqgXUTkL5cwkHk+uYQ0Rh9dqovp0WwwQFpRV41Upnt49XJhqg1VDY21D/rLz5ugv
OOAD9R2uMMJMKAQAu2xO6lSlt+sGt2hY8v0IWEfAEHtCqYv2KpFzOeYpXA6wDTLD/GkJnDZogtar
nbsfppBDPhHFhC/K8f6nFzfawHHPC1c6xZe8O0JOA8URv4jXnJ8YlIZxeE/tQnn5Oml8sSF5aZjL
BWsvV5HJiTT76z4mf/Zi/RRyvD63hEnpcdEsDzlr7xdMUA5yl9DL7O4JqKH9AoL9037BT2jAxSWm
xxRYMWsJbaiHoPmZLDv+G0DRcNLjmoS6IRdJ/Z3t9iChNJHza6MTHCkyz4Yt1jSw8k0lPtD94DCv
N/rAt8dX1RpZf09eFyCtHGnxStaqJ3Mwcy059la6t2Me75jltiB6AlYNLZPdukVf/RMsfyTfkd5/
uTEjsn4ujiGScKDIIEMGbGRQPrHaVkJrMd9RRe4qribsX+2lwYS0Puj6ODk/6pykt0z/W99ZdjKv
P5Vvji020EwZrMxfeR3cubWh0E/dLNNHIJVbEkR3YAyetUNCWJmx9bc3Euc5ankEhHzsd0frp4Hh
ZcnoV5mI9xSrGuuZiuSId6qv82yPqhGW9K/51+K9+UMELusYmP9dwXUm3+cfthng4G+h0cSYnGAm
X0xqt8Sl1dxoFGvqXrx5D57IcdUh6neNIKZSL4vmu4Y+9WX1dpcsfVI1e6VCBtDytpVFeKDkluj+
C/hc+tJ1a+qr461iIbBBFIFuGsXhRMtIYnfxk43dTs/V0nFOlJGKM1F4Bmirp+IFzolAPB+58gir
RR/6/ux8Xy9L82HZ/wpCin1f++c64urBu/1m/7vkERCr+2YNoqxXshM6M8/KP9nWPLTN+0j2H/Fl
zjPXLA1LA+dsWf36c6+0Uf4ZJzJ2EJ2Lk6VMdc4plH4WIAYpNhOG45ogoEGYdaRyFydPjd3rSbFR
viiVkZFXyzFcFwmevgMTM0mlNwHDjsIxPINv7Kk/pik4SkyiMh9fiy08pj6drL0werlchP2ztK4m
axjwup858siHeDZ/rEfsWzXSpd1th+AtTyxdJNuD4jzC1BlvnYGYuSGjC9tMD+7rLQFUQn23gSc4
+lVzkVX+IdEY7r+Ud6XUyvqm8KaBgpI6O059YW55bq50Eg9bSrcXyLl1aaHyKIMMKm3gsleV2jSk
2eMJyfBXR0AULNOlIaV5yUw1m3AjMWiMA8oV9qg9+sMti5+DGYbAtfeJLhoN/yKQvy7RyAnxOQYO
LHSKN9iqEqtWG6BbqSR4IQJ/nuFk/OfP+sQ2NDRpqSi0y02di/pblOmQyBoq7dIRc7Rl1uStt+LT
HXUA2D61QGdKUko7q6a+nsmN9A8FdaCvuzLq7xzUeZ6sXBY07TLvY7i9hynLjQdcWiCJhLBtPjII
rty42O5d4TOA/XCcLSqgOI+ksmEHFiBoMWxHH8SC9dMVxRmn1tHLasl8nLCrzEbvd9YyOfLuwL0s
+dKvuAjMFOMpNJzUEC42SXN8P/iFMbcoVN26egXhrlpz+XJONTMa7WuL84H25yjvHg/Z8FNdZZGu
ugAhmjQqRDivbn5ZxYT0VJANzS+PvQ9qbM4dfYT5avLBjjsiw+uPJTw7rSsUcynKW5KZpSuqz8zv
sK3rH/MXgquf9EBWnNikcoafibNa4GkMTqPh6TWR3C9JxnMfH/y/VWRNieNJ0nU+FfJ3WbWmC4py
pVB3FoUQ8BOs+HAbX+p+rvTM+MAgT58waQlfdFCcWnViedzIdBXhUwmI810uh5kJaHMfZtFWn5Ex
kOqcssV9UdvSD7kCxnps3ctxk1tKwLYtugUNhAwLmW6lR37ViKMJPCj6s77s80h4CanO6nTAve8Q
75qASTqE8vVeft0DuPQG5+Md5AykIcSUkKCQhPv9wbAL1Ln/iDZ8v6OskIugIsI1SgozEeksL+Me
1hokMiFIJ/CYSyX9nnRrkwoS37KoKStyWg4sPgTMX74xi7gtKnjVNm1+wOtQlcFkbWUD5Ggrh4TX
CFA7KwsqMTZ1KML7zM3tOFR6gpHP5KjFynWx4mP0iQavf4PILrnL9yWeekesOoLWT/1SwEUfJVGa
m+7sUECfzKTGxAsCm3no1e+d7bfOM6lNN6ah018X5CiM1gqFQeKsETZ6DN1lGgqwkjLZKL/8Jqbi
HhE+nrEfaTlNCu87UsMZiWQaG0W4D4TpN9I8m/trrggRqyzXvUS+6ARYjKWFm2gaF/ryUIFBaM8B
bND2/qRAyRXsVvDguxoXJ69gmH4NbD3iZD+34J/a4Q2g61l0YEp77I4SDUZCpg8pMN0sOS9yL4zV
ET5z3ppofWwoMYxT8pmKhwmzYz1fVbmurA3vQ/YlS4YaA0uiYTa+KnOn80c6Lg8e/qvUUQZajNUq
yMa/khmVpWBS/Y8Jp2wnwW9b+SH2w2XEBb9b6YN9VDcgl9N7nZ+0VZVaF9MPbbl1/egp5TF9uofA
NUtd8cmnhBQiTU1GAe3uoKP9bCS52PLTRtzxnhS5bj0rfK5F31LSBkfWGzwL1m01FhrRJi22zMd9
fvGdkolTbhi8FIzQQf76Fd4q1zjKvlXRvhjPHLodcMKP5JyHEkCT6gR2L/NIUfBizUwNzMQcCkY1
wF+xmC+ldOSbKOj12gtRkxMy5tX1kOUdnxHzAxz4ULaY/wpAx4zCvRnYXfbVJUqXBiUeByjPEcFP
O1KkiJKx4/KbJ3ZhgEff4EkFHUDvVbJgfTZ4veXYYNyJXtHwlXTQa/UFPeYQeZ5C3UdZ9SbfIzs1
cJsQTFb2o9u+SW3w7iJp98uxulCmYvgiCkU636Ya6/UwWTDizYTzNYMLulrizrVCejTUyFO0QH0W
hwusjuyCUN5gKS6uTeC85kkpIcLlYK3jgnuMUhlXU+tQKcxYj20GJiKu06fFoXazO0Qjy4LCHIka
kXG0RMV+qvbvhwxT5bOToR2WMuOLAaNgcUiBfr31NVse08jE0vrCwh14lInEOlZG5hVPkCBz+7Fj
02J9PGOCFcwPDHpbnMQMvkEm5744HiRBqbPfZNPcBuIijDaIYXzVGe06lZMaOVJ1ROONdRuPNyDP
nemgNjntrm/ck4K1VfXs6ozth/QU28qkTFQCA/2/he08vf546jmafVRibJwG2ZrRajI6bhiYzRpB
hb5a7kxLV7x4n9W8APOAZC2Srhy0d3mU3Lavt7WkB6srjgiJ533gUQd/j2rRpEdhVKfY8lSEteZk
r90mcPUmGQsROGC4Gyd4ZCEMvOzc6OmYEMo0gF4D919zkfTAwJAKfZ7YDv0FQX7w2QHcQTNQQiZc
6p4wGlmrrbSmklrKZ2zJC96qAOnax2JtW2uT6nxDcaXWxAStezqWtzrvsBwxAng2MNWM68z+n6la
6bpMaU63jSYVulhMODtfUSPZ0i5E9Ed6M8ZSgVugG0MgI12pyzTCY9sjpNWZzMwJO1Vqtj43PPSc
8fZcYycuRMTEDmBmGWTwrdKERG+4BhwPmRgvQ+jeVAB5tGkN6Eb0GneZ+L9VkPf42CEPqdCy66h6
K0YQN1lk+utqQydfVe4GZClMWJa0yLeq62uoKuQSiQ0h5N1ivSNkiGXd2RTwY9G6EZ9vAVUcxT4l
pQUNyEp+ied3xJzKrSNFK4XBi52ABD7CTn3CSXl7YJ518vwZAgGu3Bbbwmdgg29Z2QVs5FOmfW7D
OtQ+DRQclB1bcPlQTNdQOM0Ycod7DJn22q+g4Fsee107OQEIn2knmBQbSxOGUNUuiUSKAsYiprnF
MhSqptD8iCf4HK0ltlAa5+BO7MfUlFUnBgt/9p1f0EDTs7AyRUmYkC/ODU3c8F5j7iyqf7+7gpGF
M49qZSY4wNCRH0uX7popc27bPSz7MueS6COLIX20T66M0LepkC4IeF6hC7ZpnQnZ+L2A0GhPmg2m
0+1v/0SzyhkQJ4l64TBNdgp+305+B1ZOVl1biH+EzAclrdw43vVNRBZ9Wqdht3TvjMpLovArhN3Q
e6YWoghrUHQHD2GMj6V2ddS54r49CCfeRC+tDO6NoD40L1wspn5HwrG1fydCzhSxufLyGyGV29UV
/a3aGxT/jy15wKBsCxQKWsRKbf24KRICOEQNgEAgirMchDhbGUkl6//K1gkaaYKQ1az01P2Zhu5j
2jxY2YIBJswNIzq1DV/YFkzzKbrBKbNwiqHj1Ejlw2YeufMV2/XzWpQxi8wXf6C+5oIqI4V0Z3CO
pJ42JwN3UngxijVQXlnA/hGwl52PKBSmfiRMyR0FYKELdtkgUW6L8Y3nLD84r76mMNnhFc7YddHt
y3hCrO3Emb8t9gFKGglrN42/2Iye4/g05us2X64ap34aCz48K3jfqaGCNHPIsrxaTn3hkCUJ+G/9
md64Ezar5dTjrN3RoI4Kp4SfQ6FPO/cpFQw26NHtJd4XZb+WHaPC1Fjl8iptWg5v+WnF7LuF3kg5
aBWygO9ckFN4BWgcWrSGMI7JDk+CC6g5brRKSquZmU8cZG/wUIUZsfS7S54BciUttPEu+/7GfJbf
68jHCjuSR1SgIu6rGbfwn0ZNdEhOb1c60huu7tv/P8IpCagPxmYTlKC4zEuO2Beg8pT+TikJEJWQ
t5LLjTnVurLUoPvhwt+c4ik97xPGD0FIi3D/GuNdoGwC8o/Q7oY3fUV9B5Yruwy8LS8P+Klq7ZRb
9LFKotiyokzFAR9yxHbMT7y7Gnz/3PtDfnz+CsmNwHm8v10Rhtuo4qAcPmGinNdHz+LOByRlT0I8
3Gx+5Pom8Xp5cEc5knbge5Z9bvBejkOHqgMrCTXjTppOYw4G6xp1UPAwJ8MVa6oo18jc7PrC/9lE
9x5FAcNCLDK9XEfSgE3wbRxcYPC/PIVCxl5qxB1W9/pPBZCHC9RbKHK3LxfDwzrLVBpPwyi+D7EB
8Ht5XUep5z1ybtnLr5u9yTsl6KFgAU5FWhN9NN6rO7qQR+6t5C56vkyM7usiSQOCMkSB3AKrEoRy
yUOabq7R7SNkIQGq6A6nC7vPhKhUOZrI/4vQVZZSuwtI1uhdQ5W2N87kveNZZ/2YhVyrHFcKW/fJ
irl4t0O0XWqSpr6Iuq4knBKclVt/7VTglnngy4Q6CohlAxjGtLP1cNmT5xSkyMcEFo2MTXcFyRYi
m6jCj1c+8JTQUAVN6UJivBd2fA/WKpm3bm3HLjQnvLuqCZjN1ODN1j4B20dy6osCIPEO2ysOO1jt
uM489W4yR2nIPig41ulTvJsBUkA+MzjXT6hefcG9/+Pm+9ZBaH3rQv6csyr/TlWCHcWzj/cbHDp7
GpL03ldLLDurkG+PF+1xoqp/18ulpaIE0beFr7nexjHKkLzw9VBvP5o3HxEtMClgzJic9+tpBjX3
a1tdjO+57cX9Lkqhu5vJasWH1tKzUqk3KrlZiAqATvB06EhgVa1WG1W0W1aYwH7vdobrZMzpll8P
kFHPgFcfWTV7P9fzs9s0+1zAlSaCzJ/r3YZwGn8OPGrCtIWWUY87lj2oLpWpGEoPnd9gSZqXPbSX
9VLe6igx5Cv62qrqLneCdHfGfO+FrhahoIrKfeTPHz2jyWqqRQUhd7tN5S36TVxNiIt5Jv44GwXs
HTj9lY26ipIOrmBBfk6ZY9jYqGdCD+03cSjP7Wogwcq2EXBIDIUx3f9EKUc9SQkchQ3X+V6CWRz0
+MSxDxwlIT+orA3bdvK1iyGOCEvwjsS/qkfMcwjbD3OJ7A76UhRPt3HGbFh71qXspnBKNcnvTXm5
B+OELEryu/2IgcRylDxJdstipiE/TsPtJF8Cl2JPNk0maef1eEid2LASTjv50t+CFdeIzXjqYeJL
qtGk7ufH6CleIeEWVcmjeTfatoTaKuLxGPyXc3Bs4E4K0HYaXPT6Ge1noJBYTTM1vwo8s9iooyIv
CjQ+AoInAj+Zdvqnze9LrNr9eshqIZ2JNTUk6FwjhblW3wdA6FpLOZww9VMc2dPMnTnCbsp6na4b
rc85G826au6eKS6be1Qzq4dn3fK+146DEpgK0A0kYhPnVWx2ZSWgmdy6foqsAwMoHSx0cFglcbpm
alcow81DltZqqtgG7I2vhGSXxpu4ODX0KfeveCzeubb5T9/WmIGjXKFpDwWsEOQE4kSx01FVgDVa
eLbCauJMsGofi0ftMiBeeOgw3OUuYW/3FYP8rPtYKG5EiZ80zEQShwnQxctFkUeYekTat7LcexYQ
s2aPJ19RX9Tf7YO9fO+a4Wjp5+7rrrTvvyzzdFt7/hCzKVwnk5SS/AJF0Mt2vjfYV3zJQzJFa3NY
/0irF+TKup2j+WXCDV/t0gwuGi6UqOuMIaAw2rtMKyI/09Y5vl8eokXHpwFxtFc5DcOaFooPEgX6
+XXz+8/XG1nRc/85/Vm88x0KcFjrpQ9IqtfYep37OCrhwcKETgEFM552oyFn0qynL01l7cAbIPz2
A3WBgsLE0l6jDsyhfq1IoCs0cdWAqhjRtyKD4OZlocugQLVB6N4EzV3aOLczekp/gSOVzHLfoSZG
Suqx06lCE8JTVaOSUBvmIkyePYFxSbchsYr8XkrRdoz5mGW+tzvmnemeXh+HLuiB0wZXTSCkbmP3
bASXi0qZf0VEOwc5HHdFrzREacxA4SMz9O10uiDyu9kDH0kcmqgT7/2aN5LPUwb3vrK+ecR8vG75
Yrdl0rbuCRQs7Czqc+8tVnLWYNC/ql/Ek+8rkIn7ZqYHj5d0weQ082FBu2nVfu37xm9Rf0DqbtHt
Hb3zkwEwPH4a4Gp4L4QMxVtz6MXi03TtDWF2XGhNGVnzsuHI7Ez9D1OqSLRXCsQX4BX2XnuIAZEv
i8C/1i6kR1rOSHvH9z8qxYvqu/U6PYR8b3j9nMDkDcnc2/+AzLZAjpgsRRvexYBA/HZKJ7iX/GnN
pY3dTWZV4wEnGGBREXVrig+c8B36Te3vTc3yLrHAzZzxsWoAuSTDEk3MrVMjZUwzSYZsn+n61kjf
ETF+kEzEUudgklTasjpNTQe691xp+HNYMLQgTaR3pnTCMcobEnsrj48c9zXzsvSvfTv+MNzwZk0L
2JWGBFPh4BZNNRgQYY1GHy8c60XpkBqv0vN/KS4BKSfT0FraFtlQ4sRpbSAI6PdIudC7IDY95vIZ
6KT0hJOe1Mg5Q9Px/ovhnLOWBOUIZGX0kxiHEf7McADOMoiaGduX1Lch/QiGi6xlkrkYnPf2H0aV
M/IDziKQvlvQTah92B6YJ41UiA0z5Ngyloa176Cm49uUEuKrVNG9Hb9+h7n/NMuv6bQ1KuDgzo6F
DTZnESrTOETLZybVRauCmAh3Flo2ndPHw9p727OTboncm0XGd2nuiTb6N1R8vpK7ARBX1ib4UKkl
PXzm1CpEZ50c7GWJG3K+L0Iw/1ufx+LlnjhYROrbW+kwh48SQ8OU4XoX5K8PvZg+97lni1vfjfqS
fmX+m2i93y1Nt/jw5bEm/zCE0Kuyf9wORsbvttuEpxCOaAKv1O7EGbWKsQDP7pnwCJoaGaI1Jzxf
NXaIAIwXggczUl2sFD/80yTOaAkGb6na0eBDkYvxBdvaiciOlF5+KsFH1gq6R9fmbH5tj2+Kcngo
aF+03am4Y1SReBVUOtJ1vJac3R6jVo6u07pYkZNCBjGZLD+D8eRxsI/UchF9EsBBdKAU5FkUFF+m
pk2HS7xYwxhr37e19HblZrU1ngmUKBKMYtkltWE5JNGEXhPbmsz9k0X9pFR3hfasKwz23alhBGxH
kNv4t0I403Sh/1q0J3zrVcX8mz901F6XPkDPtyER7Q08hwbIjeIaddL0u28pO5+OsX97AEIhByD1
2CGDPIfP3ZQpEJvB2ESmFtWEzIvasU+E+zvn7PU+iSZvpGR8YL/74zt3YDIwyEdC35C0mM7OM+lt
sLP6VxiDMy/IeUnZWGfLsBOcRJ3biu7m9Ct2DFfrfIlgaL5PjAIwtLIBDmxTvsMh9YOeTZtlm/4y
v/wvXdqU/kTcaKz3WGDhxRTX+0Obbq7S/82K1oMjrATvf1PWiGWACigQp+pFxWWBVgdg8fYg4gan
zEd+lv5cdtQAezhJrg+ARS9dgksjwMEUUKk5gvvsG/UnNqxJQz4ma51Xm0M45SMJ8lK5iD6F08z0
WPmuLNd1NnB0GUNfgtp1EuyKAe24kIPMlJumXmnpUrHk9jTOmcZZ1UY+A1JNCrGc3/Q8o8JAUnQS
r+ElLBkBgSVjC0UcLl9AAR4y4SFj7Qfmay3fSi6Ziewt0JncukTOhCHErhaDjvelFUsSs/M901tM
mYUrWrLdYovE3YatwlHU761rOogaeq3pVZYZ8QpSyxQPbkkweeSlBRttvgImy1wCo8kINaW5psDX
XMSHdeyxxPVwZRzzvE4zUfPmJ2XEJAKQ8Xt4ym584FPKbbeQ/cVthE46+5fibTrotBFiSKvVXsiE
oyXjzLfFXct1d4s5rQkOYbKcQGdOd5X+l9XO24pmCJ/soJPQemcWXGCMe5qA8A2oqPEVOymYxcMT
/psiUCdGt+KjXpKazBLRv92HIMB5ygJYad+7HKleCBOxYFMnRpx7RXVVBxJbqSe6XARPg93SMwQA
QeTC/Vt9bIpDvyH4/Toy07XRywNYCUDSTEe3Iru7JaubGp5fQtkmmaA03USw5wf7exMvZ/D87mQ+
D2Knr7buUPwKE3mMxSjT7ccHpF6H7npqIjj9dV26KhB4h9f8eL1YtU5v2BwQmFTC7zDUnduuslXQ
JBT0BolBTH7fHQHFdYhxMyHSAh2+M6kjmWW3Jkh6X9Em4mGkWPjyuxyc5cHQPvW7RXijQx/xx/1Q
ZSapx+UZmu0EOvvUeHpBeX7A9iSnR9rP4Sj0JcdNElxQMmkcY5sbMKEt5zPz7MVXe45/Yo/DDVgP
AgEakqwj9+8dYRin0INWRgcnbFLT9BL5YEjj4ctrBDxY/LSPYRo3PC95tqc58aa58F7xdx3MUbAA
EMrzr0gncbNSP6l24upJFPz6Hufan46YbH15pWCRDtQWE0uNHtvOSnq2hlxRVb5pqgrTcfcJfIy3
ZW6jWnJVGAR0mScLEQVv21WBhahRhaYQU0IbvorBnLk5qOgoZQ/4+LeZ8LvRTBEkeZuB30VFi6Ia
C792YBZ41gW3hpm6VHJDX2wNCLtEfcsEofIDheF4ZRyKDGqXbCEKJRkSKBPJq4lDO4TYsezttSHr
CfveWMmfcmylj3xflFcnDdaWLXxmsFizGbUExwafs/az9dtlhLbYzLp1ZURMgYTC3tVuVoRujtD6
0L9K7eV1PlKx/3MwiDsdWTO6FlvCnDkXu6abvfPoyvyafTPUHVDTJX6Scu6sKUsSxlGq26kABMJf
dfngsEFD/cjKQ4iV0mHovxP+Ide1PytjisuKbsU1g74Cj1KAf9OexODz9ifo4mfx/mrdo9jpaEkD
5JrZ3d/GE3X1f7hGZDNdjScexFDgol+vELqtqNyTYAb9WMH3L0teWW7+Pm2SEOAnXBNNTTsV507R
pkPkt+/jlwCmI3XUz2qrbnrapBqRI7O+QzBBTYFz+hPQo20A15q56ctdkGQM9WdjAMtM3FkEUjEy
Ltvx/0JQn7GSRgPVYOPrnRh/7UpXrZaeLFIQiKZLtohSrl4qQqrGOZrsiNoEvG3kueiX02CZWUuW
C9eL2Mzq4LMwIPqjRQTJkrAHZeXd+0M+8VYntWWyc56rYVzU4Etoiz3k6+w8tINU8kEFM0H+ejLm
kO8LUEg6qMOx9zQimuVxwyEz9DpEu1phnSopDL76EcOIRr8jeaR+4RSyIliYu2s/cAzKnKSUHoQO
zcz4xwvDmTa8XukKr4RqjGNp35ejW41ifwCSKNy8+zqJ6ENHVZMgb3THklwcMxyuUFhqUNfZgU4K
nyv5CUavB1O3KIz+Hc2AmRxl1Gq/YvDlBuI24piGWhEYNjJ4zFUg0MLUvc2epfX0GEsMTADJnyAD
taT4xGvpVVfTVjsITIW1f2dyMIKt60p9MeYN9BXU62UnSXdSIs5R0N9krHuNU0MdQEEeswln3n+A
W94klBPl57f7cdiWVg8nDLdDldaGbLlnuseuYj0TvXexLE3uuYOeF2WWLDktBMnbsWwiba70Wn20
BJPLFet9O820g4/XQXAyx/ZaVE/sY3tHVowYMRifyF3XsWhZdGnD9Ynnki2IEtUdNhcvmTIKF+mA
2sy57XeSEbpaccIC8Fhfrqf24FICdvbku+cQU/TfEQPM6r1Iz2SqWQjnsTeGC4M4FhzTbRnU124R
loDJmFzu74Jhm0PctMPJqp1iXXGMoPX+A4XohUhl+aE1yVg4n3+1eGfRhe1g4NQAD46vw3O/rRvz
5SC7exKHIMc2E8YX/lH9n+kqO5J0NhX+AKeSHeshklJkOixE9yohcHE+oDxgS7XJW8ZsHAlyZ6CL
wtvrSVN4lqDlzKgQg6baq0R0320o6YG/LBNEZUG8lu+QeDnIQ8zA+PqxbgKrI+aciNo+UY5uxXUq
r09KviLFZaXFUcnnVg+ApknyyTdcdNN4nIXt7fVIZje4F7nfveJIh0yUZLd9n1oRGUR+qpmJVGHF
25OKj4dWdZzApjhuhYLz0shuTyd4DCFDeLOYXk4m2/QUtgdMaX4OAEIeqfL00jVg92j22aR308yo
N7SV1wlHviGx9UB2fOR6cK+ny05ufc59TGqAO2Q4BaLcoShgwrrUAM/SFt0RUEjhX5rQKeVkFlfd
3I+eR182v5g/H0f4SvS/2L7p4QCKdoJap4rlX5pUEjWxq0Z0MvrOSHzOBE90KFl0UjLowyeUf9VI
dD3UB3h9xkoEgH/SdB0aRTpxBeOa2Hfld+bcWvyoIO5Z9Z+Mg8hBI1XJYFoz1QWAGX2SBio1IIkY
E9lS0uAZP6Hq+q4bPba+wze6BKcFDeOalEHZfgggDfjobMNWsoAjrskT2J0o5XbE/LfqR2nb+kJf
GS6ZxJvG48UiVWpEbHWMoykR547S/02BPEJ5BARtmGe2HuQRWGNxLEatI7maferT9BWrddPQfLE2
37cNphB0KCpPokY6o53+vd2XgX/U2T7CkdNXw3oRbsUeIY6tY6psctVMiUWBCQtSude5Mh0NDWbQ
BcvpirWPVV+kgzmpz/K0ync82ZIAo7iLcO1h2GiA0XkWKL414PaFypVpuQNKaaev+/7jr/9/U6WP
IE1N1WoZcnoOXEcDVsbLGEFY5yzIHnYFkg2nMVydbpMWgNcFzMDVg74WT+1QeC87uwJ3AfdDggtg
vaRt3wobuLG3QKmjv3MgKv48wbdEcMc+aLovIFNI1d6TU10ShWUU3AlJHcMplp8RBYt5twsljI4Y
crSalYA5qA5aDMRH8l9O6MpjhhK7XNmeGoFxf+5IM2ruvDrTO9nnMKVYRf3lkP+c31/DsKwMDoRP
RQ7L6w3bK3EeSnDKx8Xy71Mn6gyg3oy65Y5wKelBDc8eoUYga4fT5ZtoKVwkKhImqvraQ8M55bSh
r28BlrKZ67/hGZqDWqdN2IIjbZIfqOhbxenMkou5EqjmaootvHCO1Sghaazmg6XxmEJ0f+MVis/Q
wXoVHvmhfO1BTqiVmPIN5XTxWtpTlzV5HEy0Q68HqJfunl7ZscjDgojfU/yLSeSOxZaViiy3ZWwC
bvUwzOAuEa72yQY799Vc6gEXNxqr01fYHAgZww562VH2BhQ9zESYZB1rUzerQGOu2tJ/Eh9VP9QK
/jLGOXDHoD1yF+oBrR9tIVeUrxFp3P5XNVosWql0fhDH7EGwzRmXHMQfs4NKswg5+Y+833I//vka
WOn9B3Aimk2QbxbcI4y+NpzbXKObt7O6JN7/OAQTqk0cRuuAwvVVpbXrR1VKxV8lJV+TgOB5eCaP
ntfBOPf3k7KEQZKcdW/yrToao//mmSfyQhNwpq1im5HzNjMOk5VHP5kZNL4fmcyaKTaMJQ9vAYXS
MVRX9lYvk2GIooJNyYubDOwsYw8fAzdiER3IkaZi2L5jPORyyq+0FEbllld59TGzpMhMqv5uWJ7c
TI/ecvopusYIqtVmg4pZ+keGoi3NXFmBJSQJz9cnd8NxLFf4D1mjR6EN1u0oumiB4+rfPckjOGZU
FJcTFcYy2/mn3jTNlI6DCMI+YWGfLDzMx9OJYdD9IgHk3Pv4Ru3hvWAeVf6Tz/2zn2L339SzMFlB
QczUVNuGzIBUgGuiAyGVYNmBNVJ3BozwoURnDgufDozwroXcWuvAlrBEcdGVfeImlp22Cmxq1UzS
8GEphgnvRUrw9aM8g/0AKApteL7QH0C4D9i/fGJKiSbM9WgmHxalh5wvQGPSHdeEvaIOOgpIv2De
BqNcuFNxwqCCEAxjGP4s3K91JOicpLMlMHgOzQtW0LwYRbCOeWMp9TMhVBPtDqzhFKHbQ4qCl0ms
0zk4uw/fUhCf81QhTo8dR2j1zzwyewLfclSSSfAQxSUEeTfXZW9vyTSkxnRtS1V9Y4nWyTzMB/CG
goVL3IxQdzQinagONRLLFE61+9M9+fg0PnvXiF0cVzKGs4Gye+8dl2npaz7J+YQ6KA1NPSElGRiT
oI6R+L7BbHz/UUhePLvCPeLqrm8oS1POJFm2cAS9Celdb3piQF5x3f/loehPdzaConEvC6nh4sb3
X/JjjA8FpXeP5cqITwTL4QnwAubJPjSIsQ9osi37D3hl/fn2uMJNhF2TWjBcyrxP3jIfDVL+GOCH
ob41LT6gB5hw0mUOUnZ0CJngkzcKNd9IybNEvTh0RqnQq395A9k9CKq1eSUJ+xwAU92SqEr4H53P
do0MhU8pF1cXs3O2ja6z2YK0vCaNwzTHlGUpVXHMknlYj+uXfr8IM2qBGewcbBIDYYnB2EUGuY7H
ZyqVa8/mogYFbjSqya+8jDnOcfZPfuRo8zJAsxrgUps+8/3gU/BPuHQ0CxJUHiCcNPoY+cjvIa7Q
q10UbQ8Yo/Bgb4srh2fwC1PfRtgRKq8Jf9I/ag3cXSKxfgY0zd2HmtoD/BLK4r5f2sPzdQx4JeCe
lHrLkGvSqbfNhiBOeOENaCjMRN5HYxEsiVfysH6j8DjsjpkXXeIBqzhH0WXKNOtS0n06LHO9ThAu
n8OS3MugRRYv/W9lB+ud9qCXOFhLcWRgu0xd1I62t/R0q33Jr71r/mr5Pv4SFJ0YaKPsTO4S+9RO
cAVga8QAW83lqUK5GhPAzIlBUjnbD+HfnlKhrFt/Psv3lUnabGI/J8euqa/M/I55wZwJklvUdrsq
mwgzGWprKp0tcRASSQbwI0s/kTKoblu9ZvRgiqka3BA6CZcv08h+Lfw2fzBTqw7RVjjuZciusW7f
YC4YKZa9cg2fNG5eUt/Gu0WKpV0RlbLeeDduEUh4gSLp7NotSU2vK9wdtPTQdYuvDHPKHXVmSwbJ
juwp4iP+guVAhPPnn9SJk4Ebtjxs7qiPFoWEkxncdV14RIqm2+l6gNST9FiCqVw+HrRt8u4q7ZaW
78uIMo/J5S1QnyY7F4232E3qhkiNjCk8aDCA1Xr7BbL1OESG9lUDQ/xVbCigLX+utoBZK2tVl57p
0iw/xjkn1EzWO8ayc9Dt25dP+HzobATFiYBzykzSr01X01dBBdKIujyR+oCVe/KaT/QbMz1z3PRJ
bB46+ThkMQgGIUVjcjg01JDaXRl+UMRT5Il7+/j9aLhHhBSkLFCybNskTrwkSozbTIY3qb0lA6Sj
YknIZqYcMY/F3mbhD9GjRsmNRTinWkThIJzY866otgCDT/jnnW3Pr9ve176BXVcsWhO6LG/P2A95
+i7K40pyL+h5Eodp6yljfEcpfbu0BYm5oTuhLi5i1vKXEL0ojT51lZrjKXmOkuTqNbFQN/t+W+AE
IAOqfHABShzr3xIT4cPR41OyH/namW7/JkLZ4iUgewPCyhKoAq2EN3hWABdjv2O666IWR8nkTu9R
2Hm0v5n4/Q4McrG6MuYgUctM98NfR0SaYBEjwUtJOYGzRi0frPuU84uu1QlSQTfzfp158qNqjdcL
pljtjvYEn1ZzaRfegAkI6jAqPzCnL7INQgdoFIDa6U/la9phIqEoyM0HTWLJOgO92Zvc2fpvOkhr
ht07gmJitGbVdgl1xA91c2ehx23JHA2vUE3JxteH7zCrNLbBfapH4h+ZPZeVek9sExMSehACMak+
MPzKCBKXZLPa7ltbb4PuMR9PYJ9XYQVbqumL+3z7aiItkPCMuJNMV+HGydZcmvlAY6OKgQts27nA
cvdGi9dIHmFXHno1md8qZaO1hyrw9aCe09lEUXw9K3URC5obP9orinEsnYJqY6RAbNSKBuwX8Y1M
irtECkLeH/ckeTB88YgRIgR07o+s92qWFxDc8Lmgs4ZKTmFL12CPR9wdpqea0gUuAKDNItQN4XSU
NbP+np2tU5RpRmA49qlrMx5JBXa5JIYWTGnAazWLIVgC9//7ewv58Y8F7dIicPIvg1j5gErJtxhe
8UhVvQJWsmFmj3oV3CQr8sNQT2Tj289UhaK8zSZ2CuaNvWhKtdM8qMdlgsiWeAIUIiwoC7ppc+21
ENIHPD5zTivhs57NiUDy5waOmVPKx2suTPy2opXmBVx7oBHqASqaLMiBzjbfhAMv7HBq+EmIFmVd
MHBXJWEWbACJq41g38aYxPKybBvlJS5PM81xtLv3SOsbCBqARZGCIRo225IfsgPw3TIptkAZ981U
uswp8acoEdhCQGQ3P7wuRIg3rAG8fX2cO5+svtgTZ5Oo9xycsbQh9s6ToQI4pJCeSsQI13tC/JOR
ETOEhdVJ3gNBZdwzwWywDL6DeaBoAMQPqpkzJ0zicyTMcC5Awer/oL5XBZ6nw8sYMCfZONjA984a
clSGgzEteurLT8GPEJqJdkSJojxAiV3cnU1OGY+MN1EDlXAgXv+O1tdB5bc93u4RfFj28HaN6R2Y
jGlGVB9SHbKK8j4IdcqddLeNN4o2qyXrR+eVs70mK6mnwlv2cZ2W4xVpJOFQyhH4HXi530vKJPqN
8mnxag9atDIteM3LPT6UrbgQbCg2TtroeL+qHcQ6/z7bw2lHVcuyrw2gLpM/tdy8r9VKjy9/H0E+
CA9jHh6sjVTOEekH8POfjcBHxqG0emZm35jj8xE2NrGPOgOBPeC7O8X6XEHOx2K6VH1A0SfP71Gf
+ZmJzDRXWRyqi7ZyE40sSGWNSRTgydNoCVnfv4oCgeEUXbNR4ej0iNQG5Gn+RtRXQxzPR+ngjesu
GbIWH5oXmABeRjaX9lx+D47f53dFRjKLp+MfnyneKdTPPRKSDrmYWF44e+mXjRBN/nYWZMUbvXs9
sVT4gXEfwpTNAvRmB23eZ1XT5yEkVrfG0J9PLX4KbXmv/9vg7G9X5mCltCW6I6/A9Yw/CyytbLaS
35AOJcFdByHw5BhJRJqZorVB/Scrdf7XEN3WE63it28PSiX+HPMh9C/yxviNB4g8IUseeMNDB6L4
fnrLM6W4YNfaK+bT8gpbpBdiM7rnZZNomjTUvdoHrt9W0VW9jfir7pwnaQv1DaXn8r/r6uipXW4P
V1YsGGkehvWbER2TjmsUB1oXIQTGEUeTYMMlBcuGzCBsn7Kdz5df+Ll4E3pttroKqFGDpPg1g/VT
AzfzbZSsdHGOzMSqtYj2s1fbiYWD+/HP9DQrB7WvrzoaMXd9X42h9G91w3LYH4eNteGeoXtoesfq
+9+gtz7jF7bt/KrabvmH15IYVvchdBXKng3jWxjP8gytfEvOzxtxpHSR8IzYEBroQGuLrMAfPwUm
wD5xiurTyObMjUZbZUrQL58Mkrt2zLP54JVeyrrAMINeHLSKhteiXabuudGwVa3pGstlJfWtk2oQ
srzcUOrXcN0KqfL4vS34oPcU6WXGr6kbGcnWsw2Y5ssIa/R/nhSKDUEb4rqnS/ljfYGXXsN44S0s
+XiBFUWXqK8knpZiqd40hKFTCwAUQNWot4K6GLx1G0yvWjLNLL+6KbcSQnqyC5vkhSAH1UuRyvg2
F9shXiXe+nDpl7YoVGE/V74QiLpaa0U2rl8MWcg9n1YPItGeRWxJe8qaxfiQnJijFuAGUUg4A8UK
HdyVI1LFhWyv1pblQyNRIzvxI94KfzqOsdOlx1UaoNT+LMdVj09lpEyCcpFlBBkV9fnBQ9/9dd6c
6IpfPuChSx2MnmSx58iuIxIFXCO+iS/b745CuH0MB0SQT6nA1eN+CBaRNeH9oBX7OvZBaXuzEdH7
IxZCfRV/IEe9J8i5hVe29NQiWzaHHM2O6727GBOuUSfzLFu2/WDFTT/e4xOFrrnoBrQ63jSpcelm
tQi722Fb0OdpFDLVLG0xzlr1IC9vh+qLJh6SH97LO9FxBNlUxTNKxGbCcaelFg0Sma/Z4R11pmj3
9YhqxDMrg+6vA8o764tGtp6W7N4sNdFzeyRWrxMeMXcmGgednqV6fqFScziIFKIcT4vpLch6u/I9
pCk/t388aoQN61iXgs9BykOF3hAvjnXt06RCw3t7G3WLkvFyYKY8xaCJE3mqpYQad+HLpNAlnonI
ThrMiUsZMbrNkwLykxrVAnQ0jlfF2k5FPdJuQ4LtescHzuGNoIteSH+UekQQvnPBq9CUS+875WCw
X1IWHfx4Zoxir+Oi40p2rqrXiDTnuvIurNfusluZwVCkT9YgsIla7k7sRjhnegRE1aGVNdFRYsUF
0Xu9ZwKiv0550uCla8TueR36IEIqSdg/5z/xTivIzzu4XKOwZpC5IgaZXa1KtQx+3Pi/ZfKiW6pz
ljH40XV9qyR+O3KGIwMbsWRNSG3umNHdQhHBr6zTg3/RkzQX3i0uFQkn+/2QgvTmbg2nmYUPXS2A
57XlfNNy5XqDaP7/Uw+tYyp0OHwtef32A920tSpubWnP8HK7g2t1ciwr9gbQUQcTZEjrmL8vl2V+
jxpOl5TOfCSUSmNTp9OoDQBRb6HhsXcX4QaINgOjvpAYv/GaQ1TkFZ3nZ856/xo4+wWQkInGN+L7
Baul1Bg6c1XWqL0Etsp1n9PSbEw8Vfe/5V1o0FWi4IbUR2F+i25oc+dW3PyZh23COnLt4n1Voes6
ZXaFKg2j+ORDtsJOZ0x5ujqd+HC2YG1mJq2UmSnurlVvFZm1lCMmlxfYzpCp9iSBfTBNr/04t+1I
mcI16EzoMx1sKZZfOw7XwPJwKC39KI9abTMsn5MFERvKaTMi6cFv1ZuQH4ayc1IshaV2TkiKY7Zg
h8BRz1CtVd6+ENO6ENE/KJP2lI9VJp3piCuPKyUcymI3LyyDP+sg4/s9oWQFtqvyiUNgdJLv0Cf7
O2PigaSrSVRPpseUc+Oas8T4VtvPW1ZSMWiLfyEM5ah2dM//5eo+iAcSVfYECf+wTvOG7dwe/id6
n2Ht7K1R5Au6MhWY3l2bqDEisoGdUlBzldTwtBTL0p1SDoeuJ9LduOnY+lXwF6Q5yNbPZsYU4lhO
6VA4Ctxi+AvQUUlUwC6JLEWv6Zt/LExadJ9snKUXChja1usTm0wR/K5Pl74dno0jHLVhluneynQr
S2QMQ5l4Sepo5anZgki5JoxAcudwUNIYroGuwXjoaA5TJvqDXRsmb1pi9UdPXHagzrzLm3TW2Uq1
D0/cHP46KeqFD4V1RpCrh0pUl+6Rp3/SgVJ8dj3yYCb2oKusCdL6XNC6uwL2fgvxfyYzSmLtmLOf
enWAsZU2sZVWc5q2zJciq45bFAiGr4ebQRSjPuWT4w2kK2RPKkMthBoHtofIVXXw2PsAqOxWq3uw
PWtyagvhdypmdXAwy6ORhQ73iyG200eFAgMVH3aND3RF11jOPxVrrulh3ABtczkgmURtRhMoxR4c
ZHZROdmI7FI0YAJ2jJdqwIGq959rkIJ4GrLLBht6582eOxwulBPsQHbuXTU8hRBd1Mc4dAQLcbr/
3XKE31h/hr06twsw5smmwFNCME4dl2y90OcYlkcQTQ09dys51rVpKiIzJIdwCrqTEXJY/twwX7B8
tojvj0Rktk6PiY4dxeKTZWO1TC8aLnZsvraLqKRpuPhcSxYiNrfbDt/s71OanUSAudlkKHdwUx45
cH+OYhrh2qX1E63ZB7U1s9o7YBeUmNmolG5jzKQ0PlgtutObBWN6sTIFPULi6OmnVU3xW6cfcklg
MlP3aAqWQRyc+QZh5fOUQe/GkPBWfp1uliM0s2BwoKD28bSorunSS7ucmMHZk2qM/+UIgkE2kVTQ
9ABUglFAxgq7+gHOhV8Ifp/xg9pQXIANt+hsYLuDJD7jAqif2XJtOLxRKkQ4z//NY3DQrbnjlsoy
1P8uUW8LmGBirkvzVJThYm9Oj0GhPLRFow2IXyFPV0g6Dk+Zk37QKO1IVlCBx+7DpVaWcaxyCOsM
7pVwXr+2ucS0TTcmE6xLwnKH9amt8yU5zMQvfr7KXglT1rBrGFqKgVb1zhFDQAmBxDyzJn22Li9V
o+PcIZBE3mIwpoIA7oSDdbmg6Sv1knpmuIJkBMPxXjy7atc0+CdO4RSDxVhREBzEpbbzlo2pR0n2
/4qqVHnU7ZcAQHDg+xBifWr+tdj6QCyvqVlG76limIODxrpR1I7CIEnnN/Lodewiq5kUi61WSRH7
3VC1tab1MwyvtVutQTr9h2vXOTYEh7/quwTuspqbWqC7DePkOf/zpsizf8Y+9Ynkdjfb+RtucYf0
0UfIJMi3sFYIslPHM5K7FoMhXn1l1+ZHGAETMccXctXRnqps/S2lOeVemiAp8aiAMNr3dc0AsJQt
lgecT93XdAUqWZHE1b/gGze/e3nl4rKl0fyPcW39J4F6anRKlf3He8nCWG5tFE/j36/vpmVFW0fV
rS1GArMqtlHr1DSXn7pKVCoP8y/9ZD9tXs3m+ggqtdhQpB39Uts0anIkvdxbVO8XORBXu3yEybY+
KKsVfvCZ2vDXOc+NcCPwuKHR8J/n0zz8/DbZ1TPNKXOImwKV1sbW4wN3bocgaJyNCC7GV1vIAwR+
yh0qXLVzKjtS63231WLYO4Jt2Pz6i01ok3CkPs7l2D6F6KRFtaC1bLa/9RrlwfQCswrtEC2UzfZK
WXL8LP2rtWm2Se3nT2U/iRdgw9Dfgr5U3pguEsZh/kMjoheLnTD3g6VS88NBD1T3ov7CG5qIdhKq
YxRllkuEIwTtUrJEWh/V1xMg+TOHStCY280YnltixVJW3cQpw8IWpF9jSgnwsjYoZ0/WKnUemIwe
CYamOx7nTL3FQavxK/in7ehFhNpTaP2UV3Z4SOrg+A5GRKlojFHjk7RoUeAywwKTPC6ao79IPKmA
Zoq00fqoPRs+bUcr4CqbMtOXdHwZuR1fbUgARvYfFzd30PfeoWoafk2yBgPSwXTnaZij6H/mI/aE
epEwOW5l5lF+15WiJBUNlYnFu0aPzITWoZ7nGJzShIt8rPhf740tImucZqOV2lmxcHLra+/39aqL
dF/isGC0AzzijMiGUYMzVDmWdKOhKItM8vDItpzpsLdEQ31dCocgJkOtw2wmrzKiwwVza72BcKQS
adiM56YCh8P2BOWFs1xQxQJRywXnEkcpdcQJlrgvByJR+zhn9SIoZbcJt8qb4YQ1KMPnpBFCohBm
CVqYeMbn8KK2eran+TnYzSxIC4MbUdWSqMyqIw/c0UICMfPi/KeasD3aqUqt/zqY3/zhinb1wFAa
rASecwt2CqI/V/+X78UAjWrJmyzg+tpGSQfSnuPDp2sm5GYePd0RaFbOooc1NCic+HY/sniJFyuI
rxhudW1p4r5i61oyliRwtgo94Z40glTkJUWjOgKstuP2ksZUlRebdVcHfGNwFUKxLyi8eD4UDJzG
qq5LYxNA7N4SZjVmEjZ09SL5iZiO/C+xZrZiHfA0qczgPfmFsxlKQrNMK9/zjnuE7Uh/2IaZw6LB
AeJYYgL0aKeDGXdFSeExGDJ09cRMjFSPEJzC5qkn5gpEJZYECGVskKlPgANz/9nNe6jjKqiHkxmq
s5hpktwfUvs7qln6mwuIwjRC1ruahWc045PDu8QlCaoLSNbGfzwviugpK60o9DdCcXO+IsWvsdz9
nRjhAFqYdlDTaIh8yjXHqHzpk6XLAFNPFpD1czuhHL+X+XpMtykEaK9pMkpK/diM7w1sgh5LRnce
aht1x+xyHbZhv7m8pPzKgHFrL8d/j4o4CsevV0re9Iw6agAO0W1oenTWClgDMbEUUUWEmzNnsfra
f1v87eoayePkpkDX6yAEfCp1Rs+t2i5yKpljYIRRbqNGj8XxI0YV7ApEKkzwSnCq8mLXKPytRvsh
EqycZ3ZGuGIRgLGlhGtH1U3dDLnYZqIj4o4vpasB27ya+qRBFySZLxUgts5W2Z8phJpRxcICuKp2
SsJXiWmdWHwEyiXCsJvRjWuMyR2zPfHGWQD3YlLZcI3u3XQACqidDz0rep6zceE5CseQuG8m9rAU
RPuNyPmUxzhwmWNDbQD5Ci6bPEkWQlDHBvV7JJ92oBXPfwmWaYBFN+O5nId0Io972gJECmnknB2r
p+cyLy2lY0Bb+zaj+e8yYO5XZf7DCaO4Kj5P1m7Hpe1P13pn2vx/U0rG3M+dVxq92Ity7eJSNSiG
2NBF9G/3Sp/GhfjXOTjMr/XMYguQrfjxvDxZrnQ5y0DkJz7wg4xWQ942yxVVEkEF7Bnlg4dYX0EI
crZxY27omCy+DZB1hlVvD9RRLtRmOx23I2N3GsIc/DozmPHRo4MzjezqDdu3BpKkEkSB98ANjtRC
pydQSdTN4WAX0r7h43pi+2iHzsj9nMkFXa3xwG+8HeuFTrNhIg2ue4jc9DzZ97LC/gntxAn69aoG
0MlrihviOnjDgmHd8SJf5xyBbJ8eBC/pFLA1QBpRbxJheQPPHcR6N+vVxawg/MahO0VGs9j65xDK
Lh+WC2clxZ9gQxCtUZLg58XxkDapA8cz99WWL7wWd0LC8f0bUqrWz5JZjJ4kuurpeoVf+ZPw1F1m
F6m3C1bsAH/rXWJSxp+Lx9se/bzo+V4iNcPcowcpIAJ/9Pl3pDlNgnt5x2mWzfA7kHjk4Ust0Nfq
vqZhy4hOLqpNCl3vTkLQ8Ml+Va3tnXe0HgDVq+0bbyU8qXYPwdX5tBaUjALSMb1E/XlJnhnSyBG8
57YsEV6dpPeVIki9Gy04gu7UtBX/iIvC66g+0IYDM2nXwwbLrJ4nZftZ4CI2MYdHsQmDIY9aUNcF
VaTOjYoa6QnPPalo+yRgx8toMFMmbsmIakdEwQ6wfGCBvqlf5P77HPo3CusdxNvxjAFJOHybhYxs
3HhJoVuTvlCu/GyiSJ0jpW8aRR3dnZWuF6nMkG0ebsnnZTf7Az3Vgz6aUittf0vlVX7D8rRlvd2U
ebgLPb9UEEeSnr0BXfMqKt4PDQ3xoR/O9v0GvcEnPFcNxkF8Uq8zvuBDA8KrDlNAkcMR+zjXlYjH
42Ohg2cTUat6MrvqJSI4nRUeKyVrsnZj6CWYVM7CBuT+dw5eRCLEvmpO9Z1UU7ZP7DOKvYVOzCxi
AKDwUYwo8nuj3OC8EV4pMyWV/lVgGeOPbJNEmcdoaDKadXpkKyTJPBBXzSUH9vmdGGDgIZb9dgGl
eIYh7M+HkoJFYUCLbZo6EBbxWz/euM/Vti96gZFsH4QVn1HhYIQiDbIMGH2XiW7HaWwlVkPb/+1l
89glFik2iLx4km9uj+iUvVMFL8HnDbRJzvtcKjhoflU6DRVI8GtjCugnGhoB16klTnh+PrArdKsu
pSymC0vAkYFvsynhFvGVlTw04Rb+KF1x1CIiuK982xiRUEH1FDxodp/8odQep1RGYeuHaV7XZBJk
aCyCdIWf2JrE1nZS9EfBjJPVirTbxubHI4OUb3a62PgpFAG9TaTE0bxDC20c+P599pXehJKopQma
8MZxno6j4srQr4Meb/8Ahs7uGhY9xf5xfYs0EOuY6kT9EMoD/ozn3Q7kxj1zoyTj8shn0YJYDhxW
v4RjSMQKPumGURGxeSJrsDg2g+/8xm7+D6qnpcAS2L4XO4fz+3EEHto65rq1Fo/XikWjSjOxfh1M
+AF5Kdpks3UTVOoL3IqQm0CeUsXZ+J7IBVNN84Mg1vwnavUK4ylqCv7tIybHbkAYiTpkDmL7cJsS
nB9yqJ+tysZNwNFqqKrf/qEsGLchVjkt2bx6LGZGRkxSdtFNMqtHPJm1YZJnwM4DhkZqOltSnhhn
yi5VvJpoNsec7pQbXX2XnOoRBxbxjiKx986vObhT5EDK7DBavg945nBX+yxO55uG4eLr58tORPUk
00uvdVOl+0qrk7WvscDLgm9ph7uBNFrWsllRNmHjNJmPkEjcZnRo7kZZMX82DmWVUvMBC2z6wDyf
0lecrRy4bTjMP/D6SDCpTrhdZNR66reZKV1WJCdOVrWrWK2QM4UpDAKYqA3wpmfyBcop1l58YrQr
Lv5Y2F8n5F4QrhfBh82Xkot3bGuLKRW3K9Fnr701RSpfC/3Bs3r2vXRQGj70GXIz8i3pNRwMOdPw
5x+J+obAT34VzcZBhQg77rkI5UfBSTiIReRAsN0qBCgq6p4XZNQV1ji3vFecP3UfTbUu1jXAA6Mn
gsJMlFwrYdLJ4WixTDKRyQUoLjfB0SL+q9OZebm/iOuQiy8C/O/3w1MT/qP4SdpqPiv5nH5JcFfF
T2BBmlYiiUPMccXgXoeLQ/+juiIZRvcy/hHss+IidtRQ8Q0/eOnJHcfq9Lqd+OztMhiqV8xV76sP
cefnTO5anyLYY4N3whcZTe7wXRg059GgXLV/NpBWfCUhwvlsbOMPDXp+yLsl4H/D5PFeb5qhVcjn
FVJzBktQ+6RCPJB68uJZbeLTx9AS7ALDWqByV0GZ+y8aiC6o/p+T5W2krJ5/5Sjur6auaLrdCv0n
0RqENTziXlVBlrf5CuP7ip35ozYfdij4u7hoX2k4Faa3SrS0S+ESAsR3EANfFw2eC5X5v9s9taxx
qfBNsLiEwFH+3sC1fl1sFDBAzklYRQXHUmZwWdPsf3Qa+QnDqIFMUvJv9r1KGyoaM2K+6jkwX3kI
jHylOKa5VlPAI5XSgJQBOxvjTmhNaSiejEb23b/e1DvYQj/pFqE3PkMXVJ/gQjzxsI3XRTW52Jnr
3RaBZ1CSOom1uRzRD0YtFT4z+5pFZdXPyQJgQyyoBXEDBWmVOtygZCjjogXeUvy7ET/Ou3vq+p5z
bJTIb3a52Hy7Fm2fIRdVZTp2bjs28rwbyLcV8wFZSMIOBSQo+WnoWgrkHLiiGfooIwTP3DL+VMw9
bBO+sWuqMwMjiEqWRvyhSx+6kNHcCSpHZR/fB6/WVKJpickvMLBcYY5vKptWMFO+6GjcUXaqnLUW
IMdQBXAmMhki/AK+z5YCNUe9xsyYhsXYFwr43lqXfUWX8p0Qt27yQ+vfNv4k5VrdJcHjaW+8ctSa
OQW1e3b9n3SQpUnxSbOIezBvjckpY0sdbL2iTr+YXED4TZEQ7NIuG64FtsGs5Bc3XgeaIfNITz3M
JgehwusGKcBSyG/AYf9wgzlfvltzJJwM9uaSp3Cu1WVhmFjVt7WHwHumh18bO59AMw9RaI3U/cpR
ZTevoH3NFAOdH56/g+rHYMTF3wgtcZUUB0d/ZTvFud7mWhEh3VkuarbBOCoLFvpcFmDL6if/1PQ4
exN5ZtbQ5uRlwGVUBVPqQHRLIS7sna6QC2zrgCtIeJOsCY1Dq+clECFIL4EdeL5hmt4ULr9ZFsHb
YYllDQIRorteMIhqFhBaqheTir8jt2LtV+Gt6L19iDiO4pHpk8iowVRJD5+N0noUTvVaNGEpjipR
kMR8n4E//fEUD4eQBnYzn/J3plyC4gIjuPKh039lL42ODgc5tbfceBHM2VmZ/0uFmQzph6LASzyb
1GCIz6LDp3DOlZAI9N62USwcfLClltcIodRnWuRIhNC2fmLHPxoNJgE7ryNyPk9pfPMNTSmO31ol
C5AkVD7veSY+WuJIaYsP2rkvEQP6Zfu0iSifKE21LOtUL3iBRKAmE16BY1Bsj/MIVQ+ec/61wRlU
rEqiMYeKNJNdHdddMbapuy3DGuMgS+PPJ6PBfEkF7xRrZkGN4FZJasoQTLMJ4BM3wErXatoPJsp8
GUN9Ktvj+V2WMX4BH2YQlUQ+KxNk0Du7NZUb8SbkShZoACcOucfKLVI2MjT5HVLI/mHXU0XPbCF/
SzUrQsoov7PTjBFZKAqUZLnfn6MX34v3GCdMqr5+lM/HVPV+pX3xxBTapAviBvd5edH6sWZ0m2xd
5Ejn+JjgfXr1ahILUYsczv0bjuHtCXm3Lbu1z5eB6zKtkCRCjVFSfmWYAiWG3PHkgg7iFXMSyzQT
YSfv5e7nazpR3oEN7EMsvUpaKuchKMNKf2iDaR71mUVFGT8GnuZEEV1QA+wsC3gf/MGmFixD0hj0
i3rXG+pBPUCzqeVyQIupLgrztkJB1MFs1vewlg2r31rFNkQEnkz7nBCRg9Pn4hcfQqAWHK5brwuf
a8aIUfzYjnUU7aL+Llek9wE5oHrcdrMA0nagVw3+HDEcImj30vuZi8C3SKVhow5D7SRwV9PV7IlS
YwBpmg283AwpHS8oCMQYpfTqt9GERoYdDhalbmY1hiImUe88Jdl3akOI7WUr57Pb34fmp72l5mjm
QYQMUajrgPjMMZ+a1+F1h+ydnOx3VmY5ureGFYYveKjxkPfNwlWIXNIkk3BoMD5nzXtE7d0FDuWy
RDcd7nMwVWzyev1cNFLZulJua6bZcouI5hiABzk9okofuJBQoz4CM5lDTmIFP5OIsCuKveybYSgh
Yp5RNA922lsd/6+Y0AQ7XOxSdUZ2VROLzARfHyHw4bHh/RwqznQnUZRFFEvK9OquPmlPdPYu51SK
1sVC9lQ0f7RhZ9UwhCx74AylVsYnk1BFIaSnxnfUtquVsyOINNeoMpmfhYSnpq1Xu3ftbc/4GHdy
r51OFV/EufPP5vqNqHPcVKmsfzlCHAB/fKKldyTo0YeowRcyC9HILCSJSUTZBw2CYC/Mb4Oo/eLS
jlqDkilBMbBHDGTqu7XtrDcuqkzYx3MF4fyRa4I/0AmV9vjJKowcM8PEhro7BCH+LJeKiYd68rah
2qMG0REu2e+bDRcEJapX8oUAgqy3Nrm7EeroSfzUQx0S5uGqfUH4n7VBQ9XKBomc6ONRvWjuTcW8
6dos1blje3Qd3BvyXJyzKAgfCUXovl5dsy4ELZ+dxZC1579KHDh4CEeeMd9lpmTHUfYiqLchacd7
8/TEesS9PKZuBozg/dGmi7Ad6KGeOpoUsLN/z9EAi9xhvOdAX06f8JFs6+sP5G4heDihATGjdyaK
H0TVjYkfkIrovYyejp+6hBQk+ook2YHw25giu+QQ64COVqQGlOhHLFMxFrngTCLyAH6pnKlHQsYS
6vB7AYwhfhv/2Wf31ZWl2xsu8seQtRxTyAI7od0/GkYSELtEU+dep6xSz6HgsTsAzpoMZAAwdtZ7
zFetj/cyuV6Uc3j51VsljpaUhrsDOgXAfq+OZVdrI/slnW/q8dILbhrodfFkkFTiG8fI+qqyGF7D
2Px9dzl0YNiDJTglVco2uVOBnZGhkHcNq8eEyzm6IalbrJU55LtflnBR6NRjgQg12MiNnEDEQwzr
+C3HdLieRPWf/DJlRZjHTWgCt9uo8eVP1prBKznU4VLSjXKUvlFpp8TYs34P/S9TDRUWwzcRpPgg
UjuowWwTEVPbTNLP/t4bMFjOBpsbYEiEC2HBgFpl0j/rXnLvFE4ncDEytqbkmaQmNZ3aUM94D6Ny
bJ0pYvP8owCmqTGc4+pwOjmhHNnAHnnhxLHRSvQGD1wp7knWAIguyOkDLQBORosplX7z5oi1Ni0L
qL6x73xcLMT45Mp9OOeWMTQdjZ2D3vFfwqHdJuxgtS3eAYtfpfqg9sEXRTwniRPR/yF4i48/FBJX
vDtwGrw6mrYbQhbcpjb8L4EYI53WEMSdweBjO+vvcNu6GF7e1Bn6ojGWdPaK3/QBNJHVYYaodpVg
8seLUzfyxI47QkeR73PJlW+EDnaF5PvJAHPYsX4nbi4S8C384cHXhG+1ousl5urx9liju0f7WAbH
gPkL1vCgrhAlvQ7UB21LGWk/Av+YTy1vLbrlEu1PXCVap6JyZlF4i437wWEVQikDVIjNRY2xwKTr
gLyfwzWxyn7nRHSChrLri9hGhBr3zRYkKIVc0/fbpdJkpDoXs1pAV8hJikKcP3KuteJuGHtkz0vE
+4/ry49QNVsRQ02rvfek1I2Y/FeIAF7BPzVFZgfly6H9SOEUpNp4+gGSBoXYzbBsHqkLUvYx11FP
KqRxx2QpIANdq82+E/+xmEvXK1/L1gDdj6+9OplSRufNCBdlMJt/EfcZ5X3WPu8U3Bm6TFEAPwwP
WCcczlNnre4EOliGvawFiVMKuzFlz3uBWQEv20Ynh1qREJqYZENwjFJSzfguqs+oVSaSjsk93C0O
Vw1bURok3wJvBNtv3DfOqAke0CFlclLJ641nW1b8JDNVac4uZZ2EOAKiGBvyeJ9yGniSA/32JphN
N9QTbiY8weT51UDsLD69z050PxWOQMQffitaDzCupJiSkoi4R1FHQt6YwHsXkkV4VMgu82lgDUPm
U7f1hE0oSL7J9J9BmzPpB2jR+XBVJBZjRxfqGxMRkHqMCRsLitnxxojeVarNhdk0zYpAWM0mRDtN
l9U85xsAhJna4q6JZxQC2wpzEfE0sGXJowPJM3sew4dyIG5Vm9fVv6VUyXet/60xbNCP42zR5zM5
3kwPQDqDGw9n9Qnv9IXauYIdzFxw7BvoyNPnJmVS6dhuyrhT1JqvjwLCSgdCUHmkKx5ccnTVQiXk
rturBpJa8aqz/1KNSVz4KEU438Qm3UyQU0Wn0Ehs6Jff61++64w1rD7gq4STOYb+hAa45ND9bfDT
qTc6fObnj9ISkmmD7oNPwRuwrMf9PJG7dtP62IE2FAvzoyVPxlL8BjYun8XD+7ls4H3aNDzrtm9W
N1mMxdPXVowEiLUXgXlj1B6zvrGrtQCTmY+25bd9GFVVvbcS/cxmEhDiwyQuajNR884E6DMHVJDQ
DlNslJ0T5oL0x/9Xl2Wmwq6KfmFqrVfqYppwgzNJVK3TZI50Zm28XZuNQW9eBXELou/kml6nQxvV
nuy6T9Y6aJ1WYmnLdiBdNu9VucBzDqJW5Dgj7phb36skNljPudx4OjYOM6Nfxvn1b37fLvgC49SJ
loHrW4f2o7rYbUQQ64v47LU5RrRlpwYAZp6j53OHiw30Tijfnm6Yreqe2UifDHL0K7Ep4WEVDW1z
ek0d91x1omDwEOYLBYBMRVStI9ifhbnjaYRzrbqm7a4L3aSsjZsOuGtrM0S16J8i32iKFffgJidC
rbyQ2BfERNCOQX6dsSrw+qURkSU/x7BlQ8+hHsekRYUaUtIgHW1yXJ+FDHR7eASUCcdiGHMkGNoc
AjM+B0amEUWBllg8+KU4kT3yyCtIE5Wp//enEhnB1E9+Vu8hp6sP3TQMkW25cY+/z7Z1Pu5ehx45
lIYoDvEoFrScakA/jpM0eMwBEXFBocakdArQ0AQ9rpHZt52a/UCiOaWsF4zNTRj8DfCLVYxgj49r
vJGnFcKRrN/oCMrVilw4+SqoXlVPe5YDpTBE6xxqd1PBcF3oyvQO7Ci6oHE9D2sOfrSv3R254ukW
nyBJ1YAsYKI6v7Ljtl5GcC+pMdbldIlRNLZJvEQPUd6Rdrix77p6ujP43H39ycS6au/kKkloqbNb
LPM/w/wmpn/hamT05yMlPJqe1fYpTZiFghJLHa9jjObkT1zO7uHpT0fVQs01X2K/J11i9T9OhAiC
UUOak6rio4ZKOlLdwxHGy1dIsmswFDQ+nENMHmdLT4HhIuEUQonRxMC7Ffq8U8T5NCCDESP8sLov
QzqGk6HjO+a6/5JCDFUpBsXoN8xP3WeT57PWHs8zxVAb5nMm8Xoe4x5uKWkUpjuzOO/+So2c/9+h
4qaXA8eKca3scGY4GHDDkvheonHwXLHW8s2Pn5fuc2YnojHUunQkQidlZHgTICaX0qImrU2WT0Y9
Y5qgWh8jXqsVZ2lHeMdY7jTCMfQOHbyP5wBgyhx8Td9GteyepKMse1QGSBZ7GUG8iiWYHJH/rw2s
8JT0E/vJrIXhaKaAuULSohKg385xDMBqlpa41L0sAEIcHPBGUpu1jSd6DJouNvAXf+BTkk6MgBvQ
CIgPiITgsIjbZOtfgmBV0ZrKFs2wZxSgUxmaW+pWDGTbkTieFzAG7UDn+xtsuftDkzfI/i5vcX36
fqFpkXDNQCtU3TrhHdlFEaP4Ma9s+rCK0v4l5PhlofCkUL7IUXTEYSPga5jEmUWXgY/CHUn7sM7C
UBUjrwBK6PHFKO73K/CJIYWxw3JrIDgwnX+xM88yEGQ73jotCeGGFgO+t5qbVj23FoEJpY+HXjua
QGw31Zy//fiDmidUazIakHMS5qc8ySv0LvigM/h2DCOrYiYe6CPU3ezlS+zRBTTzvk9adJsGgZ1w
VK6jrw7aOv76UFzrtS3TDWc2HiESbFxl3yKVMYi69xVVg8X/rSQ5EHoZRlW/6b+9adAM2JiNa5rj
j1M8TUsPtXm1D/qUcBmUWuJ7AqkePD6US7zFMoIn8XfynLi97QjmCsz/PFKMwkBizNeIJfFd2CI3
zfwGeSSEvYSUyEjRnr98dDo5itm8znv/4hRfY1W4TRIwH/4/yAS+xlcJ4Cq25EgLlbCgIas2krH0
bNOkthobtBnN9MnT6vf7EVM3t2b9GZaXnnuScxJ0wn1UN39cih+VHmCDmJMeuSJMPcdZ6BOqfrqt
MrYrJjHd1EL9U8vhrgt2vqCOZW4DfxgItyUw+D9tSRjzw+E0ex+oyx8OCMyRPGAE4/8DLNY1shOQ
7fWKUx3mPdtJpj5Re73Cs7m1D+6lT3ppwcd4RBTLWMaGXaiP2pueqBEjjdIscexLYOP+Ph9jT7Du
A4Vvk+fnT8ke8TD9iH3sHCwj1AS34KsAjP58jVvO3wquRYk6zRq8BsFF3OuFuOvvtBmco15X96g+
EkVu+AigtMINkaiLCXFkZpVpJJcA7c13cRmBD8j+vj50XamO9TNzQBzsWpeXFumt6O7AQu4nROgy
cqND5LFnrimt2BsRYxfl+Izsl5gRh25aFStmnEVpDdGkrgDxSng3mUQW/XepG9dK4JrBwqlcq8Xy
bU61lamSTEB8fwB75d3tlDB9JksJ7If9McvOFqeFtVRBXIBuy1/OmByokNwTbBZvzxgzd9whJssj
czViMP/FpJqs5+AoVy9yYcnCNJguxZ4Es7HoHkKugaafC8gYifuTaA50VMeJLEWmYBs9pEpKEH83
VXJ8WXB4zGGvNmjtjBC5MUTeNPpgr6DbMIx8RpoWIV5iDHHhOdTkeJULtIWDgVHx+LhpsEw7ZdRn
hiUa6p9MCHk5F1prDtmlDnSF3un1qmWKJ1MctJ2dVKo9ZPT6xFpAz0a+1BRQmO65Kv+EkI9tAqx8
UNiZqIoGP662oaMxrxLtxbOaV+Yd4L2Zyss1YO+ZtBLwmLsb9Qwy+6RT9huhDS4aZluQTKJgt80X
DVBFD2WO5QM6dlp8YJH2xH7lLO9jTrS/nJDt0IgaqZBtcsDj6OqnWAlf9QHG48MhY3NW5uXjKTZy
znM2doRs/iMK2RMeJLx8NaIek/+wycz7pf6m/1h1MSk/jjfXoTDQvXkpjqbkmsZZYd7YlSquVzpP
2fv18pJWE4KRNxv/Qe1eP6ngtRNOfIqP/Hh2JujBLY8tmGc0jGcOCbv4snOasESnbGa1VsOxUVtE
BgDo4jzPPjp64Z+0wRaKLbTOYNX5eLX6hdtjBoy6G61//aUaHn3C2Ln/3iWLv9IikwPgnIPHKWn2
/0dWotxjBIa9Zm01qL1XCEHAAtt5kGK38ImF1qUDjjORlI+lRRZNHP/gSXhj9caxfJQzNkZ3dYjk
GA2rbR7twJNvCjUTbksemK5TkZHCtAq5e26mIqpYaNcKhQpjJY0Jko0p/s6vNerJcuPVL6RRgg1z
QhB+Jc/EwqpYPU2WpkaVCJfufykzY0reYBSZj8ZOUBLvPXVfVMjjSFcaFhVfXFGk82HusBrjyrQe
Uhr845FiA7choD7TExQDlpy47qAk4ZFhXT3qqD4C/X3b/YMQYkn53YXah01EXUt9L+qxUW6uuwci
W32s2LkRK9X4pxP8ZoEoZjchgWkvA5dAir+bSPGYHyOCfr/8Z464q6T7znkyO0o+gzK5Wo+8/wij
bx75Whcu1e28lhRzPe+NfL42wAgR92d1ZwouLrPdnurjySltbdpAExbnHt/wY7KeYhszTySNxT7X
E4RmTHqmWUQRGXijQ3NOBC/U0WDiUUMBvMBGc8omKjclQJsIajkmcIYvA6ajg+dpj5bzH1aPVa8Y
ldt2vzZq3D/4lpsoShsCd1x1C2xvOw+NEjpdAoiQJ0os0MUXILKLpnuOQTAJNcEJoUjwaOqnaQ9j
RNG/7ERof08SyX3W7haqfKLNVJM6E4sPNU9KVwhboVEfoZHos2BLAhOwVRt1kKlbjDCq//LMeor/
sydfaXK2FPRAwsj8Q0us7OerwYxrxPV3U+R+P/pjL3dsIhsTrNEhu0pLYzKBiu9f/P/8zNaCl5p9
ZvXGin58NWeukQ56iHgs2gXi2125TJrceKAP/fM4wPBzElvkrDpHqaGxTuDejRwt0rcOFPkdGh5g
ufZUyRIXvDq+QHYcs3VnYjNfvp3YwjD/8x/ZOnEX+0obryiGRMV2fQCxo9L7aFGh1Zc8K3ESuKfk
k+v8l/+1asVNGDKs0uzhni74HY6NDuzLF8UvRqFdTkENZJ79DDJxSOzvC18CrLuBlR98NVemu1hf
+jTE3sWl06Iv8sAm9fBzgeitZgiaYw+ZA8QCJjnXYW/mu8PptEGkH8A4GkJCZ8R1jx79KY0H58H/
UduoEhansc6kusfecmk9XoqS649DsdshYVJ00G+Fy0N/ELAT4tY1XWnGR/GzUAAYCcfBuIwVGj30
D58SMtElBqw8LYxJKE2VqXHWepTbBbJEBz6X8f8O1YkVMlnSfqvzmVlhWGC1qpCXzLyZ7P01F+RO
1u80kjBWFrZABacrYoIA4tHE+5nOzAOwaTR+HhhwGp4EX/fJLY0jWy4lhefN5yS7TP0c08aEIMa9
3lpnxUbd3CuSjLYS9BvQ1WIzn98x3SZzUxSWJ0O+i8XTh+32sTVBElwHmUwR5WGXSs4kFMHyB30U
5cVKbKrSf05uWfYCzdWDYTJdaQz8vczjNFhz8UvFnTeMEf42s7AiCXhbNaI4vAqQJB2WymsKG+72
H+JM9r8nxRCPYV0PPlKIfKO9oFFfR44BIhesTE0cT/OCBPpkQ/652jvQFb+1t/yx9RVcFKBDuQI7
5C5nN5i7Lif3acIrY872/Uq84NRqCaKhvIr0MZX5jAjfMEzHr3qLRrqKbJBZzd0Y+BBji6b0/sXF
LlGa7n+wvH6VIoSwv0e8xiVqLHm6r3LhOXGYBOBLFN4MPMB9KMt86xO/pzovhsj0wLkX2W++0oFd
ViI39acLRHKBPa4wNnCb6y9m6CHr6sRQEYKsdpI9YStvfNt5I+jToTkBrwZljU0RWYcsCOOgnIjl
sUZ4KabraE0gvUt+MIzZLSV/YHJRyTHYmPAPcZXMhM+x3yB7yd4DAR9ei5ByG43M+cEljsw1AYrm
zZKJIlyY4dOzpROT05aVpoDBoSPjkoXRigYi9eTCgBQwHHm54RFOxthqIAqMiC8dmFs6wwAjQwGn
lS4x214DcZbzo/x2HXUj3cU0HrYBLsn+fDHiLyQsOBTNyEJ+09I9w9i4z3Sbgld2Cg4e2SmLhm8a
BvIQIH05OvuZea3UgMrLIQsKj0SVNBh+oHJ6fn4kso53+N7LgYkNy8qkn2xiKA4l8cyGJjVP6qbW
BSd9Cty49qJjcuAIavD72CpWwSFJTQkl8OyIuCsSbQYaChlzwCXCKmsODAPyNuWlIspYT34EI5gz
KNvq9dia2bHSQpCc3/fvOhpzq84YWZua9sKg/opJtb4zWNI/fh/UT/4Pm8o72qE6mozvILtmPXdp
JyG5wr9U57tkj7AJLelwcweCkDZnH7tWxdMGZgG09LSQdZOpG0T+u41zCnBFY3AU2K6Vcz95a73M
I7GwW/S7k0SJ58DQWqIkdfIAaKC0E7Hioh0HpkAMbq1/xkkc2n53xC57XB5Yyg9FjqfsSbjBrw7d
XX0VJk8DIIoFPU4fqTxqgt61G5q+VB69cUz4JDqa8LuRRoFkrDj2gup/w+ZGsQkJy78hwWeLsahS
4DHczdyRzos6V7V62rV6VFunvJsrxWUCuORM2zMY7iWruC85i8VXmVsiq++GSAoMCrJZluB/05Sd
+6vOVnA+1gCV5oAR0bl6Vfl8XqLIDrb1cjsFxhVpulrA7v9oOMo2Rmcfsgc1e4jKituLkEZUGXQ/
nkPcTCr08XiIyPaS/PafLOS1CmMSuUjiI66+wPRKQrj+2VSJrC1KySMdviF0s5LEBsrDawU/zoUG
DDfqZXnw5WOJSEbPl57dA5wzRPMXaQLf3kLXikGKJCgK4iI+UMc2VdLM6gJaom9EhiZ/UIGD+zhm
ie45tiyFqvSUJGbb23CA8ePrySwoG/3hxCh7owJLr+dDz0/twJm/U10j0RUsY97po/UMEV7AAsPw
EvjoTSDGP0sdvEm09ZGahNhBUT2cAxpuZ0pLBAssCcfXTOPCt53vWPjgCxtMz/p2yiVZlUd9moCi
7y476r4JNjTua8T13JbjOPR0UpgN2CpsGrS1vnRLhwcXVf2B2v2YwgpsAgvF9/VeIM96NybNAi3x
2rKDD6DKNew83c8gscuk+NBpYsGu+YQYgnfHegi8bPenlOkL3kSumXl/ZdTfVGS3T1Oq16gOFcoR
ojTsjj87s4QtysP1cMazHIal3gq7OiHmaYQJOqrkNldy4Nx48CcL/uYyatSJ6mf8jhR2LQlEtNDA
wTX981fmvoDRcQjn+1F1ofXL0Ls1LnlFUh27IhOi8dy/9iLA42M2xOqZmaE6tH7yDbgKMZ5I89kN
ruIMUk7lFM1djahIujbw6hQ9D2AzvvGdsjBcCftMzU8eoeRAS/PIsob77l9I5Nk8xkBhac0J66vT
KjZNHNSEN3bWmnvRgKPdE2EzCHhkLwznRJuM7lj/D/X9pSU9Bd4a+EFFDO/gVLPXa8OTNOsWmk5B
mztiaYH7G2GP9bfWDie4gbMMszCcAwhLlMj/06nXzOAjX+qqR9eZlIzWOoIueRlzcdl01byJtknD
zv+RWJM6+kw1NIO+AtOApHzNZlQcrrTz/l4tvekBm+IB4U89AWf+bInsjyP98bdXTz0mCwTSPlKJ
28R22rG1NvtMjQJORBuZHvqPq1UTNQqadwxIL4EWrQAQ5IZoK24ADZDFm98hwxdnsGR+SgoikQGA
l/EBIrsfRjza0kB9zpFMSybsIgGZRCZJ9D9RB4rbFsUP/DJVkHg2lMktFfQNFE/EFsEvdhz546M/
SJ1WLouP758vqgF5RAGmMypwHAbEH+wEPn8KG/yojg7Psvs2LX2jQ4WkbLTxq9jm+RVIjwOuMagW
kOROkbBZ+AiIb1Qk58MdyQ+Tdc2bqttLFtEGV8rLAPZP+2lrYriT1M//AlxahB1gt3AVlFY0+L9/
C+zTvCcFj2wxDZlCr6aKdqvMPGFWZJYFipi39Aie7etrJGqy45qRvLOlfxI/TcvqrfRz3b+Nnd/2
PbnhNZGFVBatiM58Zzv2oFmhzKxPzuval/Vpayq99W/tiDe097D+kdFeN+Eq+W3kWDj8sfz5tXPx
eTuBskv0mcG/nwSpjcJUWjP/2Mnl/O8ccAou1V1WeqLhP35WF8/AmVPNdbNCB+17EZ6hOEfgY9Mm
0Svh1jk4oFWPDB9duBjBvbQq87QRYqAdQFn6ofHouNm2YvaqpEoDexuNFofUgBWon1KyFzwtbYnW
Zh24XeyJsIFuBPusk8RAxj6wGRcLsHdOzmQP1ReC9MMuVLG1pLjCqbiGX39xRr667n2eCp54/RN4
3ru5dCgPjDxhb7rs/KWRa/QDmqVYv4MC0Ns6DqYHKNBtBGT9AMwQ2ng+L260FI1YrNSLtf6o+9Ys
xBinFpeurWmqeuS8Zcxk1WTfSF44MyUKv/2LbOsITiYyPA/yTmWsahSHgjeD4YMxZ+rcM/iCLMLh
w2XYLbuV6erxYj2BS9EysS0QRtzC/LdcMhgWrRQK7+swxuoFbqcDj9iJlTDUI77PFt7HCLh9heMQ
YTBELuaXW51INkLExOWpIBnH2uwaydShyMxV5O34G02j5qU2QH/kwWTV+XPiMTrgFuYLsCr4FPD9
ONFE7WQ12gfVpnvsQ+6do7G5DyPyPE8hRhNad/UkkRCaQgPmT22VlC2jMyTCzMbdWrwPKfBTnsPK
HPdbmE6zMmMFVGLjcfK+y0E+OQE/bav8ZEX4eXw1qH+GFZjLlIVU/xaAkI3nOvmloqmdeBRWq4Rd
zML3XhpMgezxDoDebwviBesG2cHfZWlBSpHv/YzlZlWZMwFNg+11x66Bvuafg0OtBkaqXW5wQ4UC
yssKYZLLX8FNi4w4Dwkk88rkFZL9Q/klUyRbdZ3BJAdVMI7RxJ91rk/U5A60NzCHsGpePHvX7wER
anggaY+HHaRSglWfYzviHh2z0UK2JqX7lyad3Q/ZijxEoUJII9K14sSi8334sn3J2wtlcufx7rNV
CHrlQ4xInR56oqqrpBaW8xYGIhVclnCa9BXR7xZ5I5jaKAPzWI0boTvYirrY4q6IQbxS+8Myh+cO
vbhjYl0S3TXFBN/hTHvcexriGgBlgbs9Sl2vzhsQOOXGiGlwVg/y35w02VTSISLL7t5FFq7TV3Cx
mn2p+untO9oIKTUSNub6Vrw47jA/Zr25HqAyPzFvht0cVm1bZhRq2jhEkmvIaGRQZZPdslVs8wgH
Fj/ezNy6r9yv7Ivd145kQAje/qWrQ1w3MTCwGOPxy2LqLZIZ1ACLlTqpda5SP3VfgrF4aodVQSup
iGJ0fQSKbFc6NVVRoPd8hDrEIRBGSmECcF/Z/YazqiV8BFiT0zz6CRSJWYV4Z1dxFxu/dggZJcMX
0VospMPZpQDoWFCXRXY/wacf0q1QCW2w6r6PXkiCRha9KNcAICDyCzZP0W96geJXxvO03whOsD8n
QtOZMv/0Yjn6n0PtKLxxERsmueTb0nsjPJJYAVJq3z1AErZ89gZ0RDcQtNKbyX+yy1eldU1AB4L2
CfEvIyf20jOl/dfhc7e4srSNhA+4NrJyMFoHpqvt9NY+Xzr2eTOYMa4DtPFp3mymo8Etgv754Dzy
gVXEMIRriFxfzTm8IFcuf5MXe6z6VmcnJYADcsq4Kp97iv30WYrpfhdf89B9WHiFeAHyzLSPIKKZ
Up+3+lM9Ia0DZOsnRfjY84996hbI7/71+IB0DNgYX1hANsoNAuQagojQB6uf54JMXUlpcrnEFOV5
HzdHx1Fd+jqQPNdE8eHTGDxzX9z5ka1aNfueTriUBlXNKQaLWcLqcfrcvVcnTbZv5njDbCdEDYFW
rQiiBgLKWFGhOnJNYNqzdHI0R638QafNRU/5a1syt2Xa9ZtjlC9dmk7GeRqsComptHDJr6Lb9N8+
zWCPhp/S7Izdf3+LTxHtmCpyIcUHe1Tt6SU+Rkc6hE+JUP3f/Uqvy69s0iyR5xhK49yRXKcBgVJe
s+2Om33HK3pCtia2Y+QdS8ZmjpFg6cCyhEUbu0WRHcx2hzQYpNceWQSP8thiGOkPSROjlU1dMvOW
MsRcvbuBOd2yirLwoLTxcjARB6iK8AtOFI4Jje3B+c0kclB5kUZoaEWSsu3Empt9pnnC5HGdKMOp
wQY2P4DhtsWw2cBgt2XOUIRoUG/mi/7HAo4Qou1hrI/F62ySuzvVAML+dIyRFFhbFh4EftvSCjCe
paocY8zimxNvYU9jkuM41SfbqTxOAD16xJcAqBqyWytF+Icp3EEwlRADbsVFJVA5CdbiLyUzxFdG
bJHxoMLvVkkYwqKrm2XDQLViuKhxFk9PmL5ql/2avQQil3T6gIiE+j5mnapSMyW6gNGFM6jp4jcM
b3+pPP7JHQPVzMnCBfstNonSuf5J1wmxS54Qj18nvtPk/e8YLQQKmdCySCdbzAAjYb385qzSsq/p
ju3oWRebF49/dnwuSm/09TE6qnKblEXxN2d/DqgrjGgypXd40zjsNnW5fynXiTR5WvfA3UyUwbMO
Lpuzf3KFd1BMNE3j2F/RHWxhxAUki9wvJtpIHTbYCySq4D8OcomHLW+yTT3kF+I/8cKwpJtvWMO3
0GfUuAQFevMVLQQ9q9oe+QQmyZJ7Y/ea0bI+snRhJbaOrggref7OQ4T+lFzzVbP6RTGsT8khTdc7
0rhqP4cmKvSdsBQiT9fqN7m1ZY5RnMWEkftHfiT2S/468HwWCP+tXl2gq/QVRvz4TLw4NqPE7h6L
/mpNCFvMoXllxlW99AWDQWcElsniIfVmhRri9Ai/rgw2Yn9CR8ZPzJdio3js0kIqcPfWp5kRgyVp
5DLxRA5O0/wcWp21ikkWzkx45R+jHZa0U6Gt1td/LWLOpPRbPdesqRH0qYoTSPMGVVHUGBsf8VhZ
EA/BFZAtuEZb38o0hq8fKj9cd6itNjNyekt79a0/zLEb2e7R6O//U7u07dEJCgsdEbf36w9mkZQy
YVYfklqQKsZgZXNdmjNWwfjYKOhXeY+/2kt5eRlTXjZsO/SbY3iM7Rq+St+ApQmyOpIUW89+x0uT
feQhwYWh/S/Ly4Zi/opDf7ssAGvY0KabcPgCUu7P0R86DERkjf9jhHwC6eA+LjrYNJGxEBcIkZue
FBDoN/xWspvjsIyIV+Tqt2stnc63lJ4eFQ5UDjdIvoNFJcB7x9R4mBRy2g/7YK9MzPJsx0J8yDuN
9Um3fdac+/QAQSfaFPL6tTaFxStC1X+HXFaFVmHVTZ65GDCdLXu+DBv3PXeOj96ZwoPmBe6yWaLz
Aq6+Qb0dppqBFT8lW7qAyiuulqQVwa/V0AJgnj6K5PrGecOVjWXaeNLPk/KSwCGpxC8uW6na12Rl
ZGMw094TyGSsKZCFIVbUueF1Q7j4XypEVGMCKr4hE+4g3aeu4pscFaWmdt39x01WEbIw5LM0DghH
ET6EeFghiSkzC/MgUJqvjNZllutrNV8Id/8aWIEf7zt+92Pn11z0DGLf9LzQrqWwb6eX1UcPqRBn
NOpVfXr4lIQY2CfNz+1XzF2ZlIZ8MkdmeBFT2n3FPHqIMrtkYNx6ieEm22GxaFnWnSxV6aJ2k/oA
B3Up4fuk8wEp86ni81KNy7U4VgoTxDj94BO8sFkOu/X22eBf7SeVwg97XZpQ1JWfnauOzgmfC/47
Y+5O/sc16JuaLjsS6fmZgin3VY14fsHsjC+vGOVCfDJMPboK9+tU5LFaU0A1y6fz3ly5JcdUEd0c
Z5lqujwJa9MrJd5wZPVrnRX7HehjGdM54zOhSrfYLpGuKyOrbO/9C83S+yesKBvsOf7kOB7FD2SC
3ISTUMH/xujieRoXFl7n1dWI1afYhrI33/bgn8530EDnJUpqF+CCzQqlBKBiRIqOKTcP9n/SDQ/P
AAUNpEB3E9MwRxbyXTN/KZSHe8sbt9greqL0qm3d35eoJlCr2H5Qz6oW1k/TPlIAofco0EjK1dL9
kMDaC3Ekpd4bp0AqLfToHg6FsRVbEiBOsJPWd1Iuun/fyCWM7lpbimYCHpjE3KP9MC/88xhwWH/J
wK6sIFn2IromN8kLR3yKxaeJXGjFFMtoNrrAR60TurQCdqgrpu+1ZzWmJ2UO3aOjGMI401TSdgBq
TtQNkDZvldX7WIUJ7UmY7hn3GGogjjfM2lMXq17Xn0K2ES9NJn6fqD8fz4S81AbKQC25LBTNLYY6
AjrO8EscSeWpv/4d+VV2t/9ZlMolB0rnLMz+jn22Kvj2rS+wLeh0aI1lEVRjFCav1zR9c4XyzWbO
CeSkBTJ27xa188ZBZ7WzqXw/kmTDUj3fq7akUId/aUnr4jSSJ41/yBYKyzE2eElAjhWL1sXPaWru
ffifcjmWV7W8v0cPI+wozfQ1SvJzVSeyD2vCBEUEOX+32avLyTNNYb+H3nxO6IFxvCvbtuu2EEWG
8sHt6UTsUNghBs9ZXhXmmLd7O2e0Q63gSe5OBVbQ+fKmIHTrT2jdj5H23sIuVcWM6owdvek10sWS
41U2nbu9zTO07U5lPRbc0OHnXpvzm2zhu1mCaHsBV78/4Dwgjxp3lgDLi/S70ljdW3ZExEBqmdKq
OoF7EZ7TpTH1XBmReCeF3aaJOEjJVLv0SE0M2wYUCU/U5Ja7CSQ05YWOLvGtVCEqMZsTe9J523K7
7+sYJSeiRTDFNV2MwDbsa1KtVHi4n5Vo7HESRk6hCVtc0zQhN6+m9+F+xQOyto22e40JOoOoHfx1
GlWIAGJU5OP0MBCklLgOXDQLU7bGQiYxpxFN0K/Rn9nqXD9TomBTXRtPU7VV+8W3p+mq+sB+bs66
fJWwvwbNxGihreerJjeIo3alK2aXj9Hv+fWwGXfQ4U7mj2BjbgzajSBdx/yrXVzv7p+U68/cEixZ
WN1nTRnlulyASwJOHvWScvkg4BHHdkmuplqF9QfeizA/mLPjPsE9/yFrg+GlxAZkYkRfavL7ahWo
c8XV+WI3sZY03s50ifzam0apbr+DBFNlAW3Ho6OdcUHNAjznpXDwFgo+ZrgB20cFkXx1qZAT6/ha
a+gQNxKOsuAMlBEZa6P+meV0ex4IXfH5pyFV/s0RSdeICZ/DMkyFoKEWyI25llCOwEtqr/ZoFvGT
BQmFwigjCuA6N8RTWl2HTcqII19y77PfialhNnV/yYN1VAZ+C82kqehLcbuf+9pz2EKO+C0p9JAd
1D9OgwcH+nhL4dM7rizECG4xotrH9l+hYNZ4oI4RSRS9j2P8LwRp1eKYl9GCR7WxZ0re60wwGKHx
GaAt3kV5QubWMQzhRHbt4RFLkmFcvf2tXE2CAAbwwE0fcduI+0d20QoV2SYkOGck+1EdwcsWZ29P
bL5cCbQUGR5uVePzxVHVBhQpZNNSOZ+jk8bqTzfRg9HP+Oswogc6N3fPJl8Z2JDDxl6CvVIrTsny
1Ol7xnTgk/bCLBjDrOBqB0rZEse9ObOxRY/IHyGnkAEMid0sFiptj+lv+CB+lGerfsNwB6ARIsgR
UbL/aWZwiimLwLeffm9Swf59D1vRTrIm2BRMONk80NEuT4TjZqLwyqbeUHakdwRMMpTDzqXeU7BR
q6v1/nuMQW6OBpXJAZqbG3AfzQPQlf8UX9lhqcX5hIdlMLU/sbz7tZOfjpkJ7j6FxZzLMWS8m9/p
Q4AotAWwZsQpm7+7yLNACcn51LJhVfjj+oxkuy4G66UX7weZtRtyeANPDqbGiZbQI8cHSKMWu/kC
EE9AK/m6dX8RYCTnujX5++wU9ARxngP6vbaPzIMOT9lkNnqyOAno9KX30LzmpIp1/94YWJT49xEJ
qgD10wmcX+lT42kRt9K5mBlYwcjrD/Ji7O9N0dC1mENH5sCrmNWPXpTdH0zerIbZxPms8DTaRCYR
Xfp8hxPsmh1uGMVSJWAG62KCJAXhWhiL/e4NATO00gJArLm6oK3awoeBsE8EtRuFiKCLZGfALxoN
7gswQlR7ce4IZ6ai5m/nchrzVNTChI8tN0f8VK7/GojsYNQ0miYlshmpyMTt+KSVz/nRcXrl+N3P
WcWjsIGYBK0V04bu0+3du+ud05p1onmjbZ68WELa6SDnOxTgTaYJM9wnT1+H0k6vxiCEBohn9ryL
5169UU5rd22O+gP6RnDZwzx2dnxoXp78wwJt42obAdmZAAKipYxfNpN6tDpnttb4bTZgFfMNn4yX
34aabReGpW5HVJxOZIyRXtL8Y4bMP3k0/OpwEDWB5FNQucYKcltS1x+BXMaRdgRKdUk25R7FtV2n
8jWH6owkYsx0i59lhAuw4NQZtmtfSlbnlQ0hRL84Jft9EX+4CIPQEiUvrCTsKbe1M73kNf6fTBQJ
OqZfrAsN6aNX6efFv5LRfzgJaWxr9J7anoy1Gbzy/G74TUSMfqECmzLGxknV/g0bRgI9Sq9KuRoJ
GBEtf4exZ4Qx0lfEYc+NH89kSGjC2WdGBZ+XjweJxuTOAKQY4kf0GA+kg8R7XdEmJ3Nhqt0tmr/D
53pdCp9oebyRk8SegQ/I1t5h6dVyFMUw+PVX23HuRnTXfKfI5fvYv98nSLQ64O+NR3b2mCsfdYfN
vNaMXWt8xRWaz5+58oGHL5Iy3F3ZNhbtw7O/a5pWjg9z7TgTPDJAV/lsZaTfzdDOci5vHbqLRMIM
cMjLvsNXWDHSyc42QLp/hYExx7MJkt6VUiofOBAmJaUFpOT+jSxDUyRwDAWBlQBVcLuhxRZHhmwt
5nPtItd/OOAU+xV9tGn7bsVmpR3jGmuEUtDdGVoj2Kyi/awV8JZw1nd5ZBwilrlgfAOceMouBo5b
mPDewlQ6QSA9p+QZQUlUn28IHHGetMj5UpgVghm+g5CDYv9YBoTahfXw3aWQ+xMa0tJdluOoVYny
48iQmkLajH1QzMl2WSR8fw1wFvJTZwv673tRcbCFS1NqPM4ZO3rxit5v5hXlY8CNa3S54PgRlY0+
mmWMulbfNuyDQzb6Lf4y6q22VvHYBdMh4ULfrcC8YngoBSVp3H4UvkTo/gtmH0icsexn3LA6SJPg
ULTR7zn4YWIpOs3EDeQZYDnOgihPOaiqxw5cGEXYmeNP72zCiWxzRJy3lUEcLTTzzED8QpxrzUbU
LHtN6cZCAqPCcKLpNyl6220/wwW+1kSjtamVz3UIkJ+6SceCTkFJDf7rmq0RqsK6mzN0KsbnLXYm
aPx5RL+FY+5G2BXkz+OoAL9BEjR119HRahZ5asJT5+6kXpc4LWyANBeoqVXYgOjqBmWsL0L/FBhN
Oa280U1HEn8vbQhtKbpRuGhy5wWKAdci/3efUPSnkd8a1PmlYCOcrav6FGAcPDatRI3YDQ6Y1+NH
QM+H3qhbDchZdwv8J4JcZK+RwTVZQ2X6tdqmv8vi/RQT1/uyw0VHhoKeuiFKl6yFO28kkH2p42Uz
nIWNk6/WYCkLBhGRgpe9EyL3nW353MNJ9uINM96w7qdEptnbo8vvUeRriOqj1QpjRnh7E6mMQ2zR
w22rxsLalSpjV/fsN9NNic89LxCKxJnmWyW3Ur77ZamzLB3cC1Efv1NEUdWXkHh8c62zYyMlq7rw
ABMwsldPe5+L0iXp5Wrk/6be5/WP5WQ/NXvVTQv/EbAeGJZjU1vliPKCA49LsNQHk9dB4W0S2qfH
ZdR3cY4txzFRTGAoMpE3Z0F1XgvmYw9/Z1g8q8qB+ZM3OX+i9k+F/jWPGQDoEKDxNZRS28lQN1BB
ZIeLelp8pHtmUpkmwh93fu2V5F4oibQqeYOm0wDjAWfkKHJ1EbRN7/1s1irkdr5cJUlVzBrItLqs
RyWgRO5YCmC286E2fg1KPf1K7/yq+PeWWfj4eL3le+EsCnX+S+xbaSdaxgNYpLxd26zA+eTXz3TA
4gdfuckKpdGN+bIbcfM++57/A8h5hhRqqB+GUtEQxDW7WNGC1UcrvqIJWzfQEmemPoEIFnfmDBlb
O0dT2JQiHPVG213SLfGPy6TtVuVq/446jlX4CyzGv61X1lKsp7ppPsjRCcL1u6oJe81v1vJMRB3s
i6pP0CW2orRx+8jUVVf9oHaxnd4SsK+B4BjItdT7UYMCoVa8CxDD6Qd6glWM457N5Qr24vH8sfs3
IJp92RmhwobXl+AKF07CoMm44YmZf+g2m2+gStYK5EimYSyAYNXSu8asUu7fkNE+YXkWc13Bdyae
213MWQjjGM+YvWzajTz8GYxNLUwQCTQ7weyjpKh2Ft+oIBTwp/ERTmEEvmrnIuRxoToS5hr6R7mt
r1oTFWjfTxxcNIckJmV0wb/8uLmDLw5TGdYc8b9QIONDecPlyggIpI7yOFnhc5TuDnPExbotxRic
7jvZ+705hNp588i7mJsvJSSyUi/uAvF1zHDbvRhK+988LK0G06ceH9lsXMkF0Ilz4IbcJgdTz8ri
u8M4x5WJkzMKzTSV4l4vG5UwQUttkJ4CzBZF47ZnP620UrDnH24N4zk2dGECQoZ9552+gwW9ovl6
vYviqGmUYG+E884GQL/DY6MabFlw/NQmQ8ZxgnagRkT//DIyxdg2W4vTFs8gzvQ+kVREDPYSHxqJ
lhiIQwo1NT5cuTar2QrlMxB5GQykVAG6WiAcGg0C9w8EkQuQAe8IKwdaYIm2KBInmtGVpbZkLPA0
Sea7sLxWctgoIscyxhRzkejuRdfA6gbHQWh6iycDsn1oMTHMP0tm5KVnWai2a4RGVWWojzvYjpAv
qTBorQaBBsaifkJKEARj9RHyZcp+2haqz3Gz6QmE6IljgIifA+Pj843Ypodh4jCJYoHdrtZgjANo
7FMlHT4XukZBnSeEv3vch3SdYEws78fsk4egmEkFcYldp6qDk3/uaz+pZ9/4rqeZo6a+QgnuV5nc
JVGPOMcB6jMRjZhfl0kdpIIszmWbVSVvTAOj8zuCiv5V/zZ+9glxoOZdCi7P0OtXUzLcfetjV+To
YTNZlqX9L2ox46sB2Eq1AMBaInyiKa2RMfqZrfEzDGMfDtu+gSIGSGEFJg70OvAGBp8jyaKg/7rJ
k1hekJDtmel2GVBWFeNVEdJ46mWpEKft6aAZFnIGxJ9VV6p9KUoLy6NDN5jVeygWPRp34Tfp2apg
G0a+iwPMzpS1N61NcG0Q/DlCwmUi1e3034L2oQVbosfQovj9kUT06aP/Cv/nZxBaXjFOKnHich/3
4hl94ewNfbtkXxTH80yz79R5O37VkVX5gz+o6ZVVa1gw8bcvrTgeNA3X5+qx8XJGqFYDAS6tzgiM
Q9Itzz9lg1mQHZE/jkKquZvb7L8RZtuwAoeVenEQ5Vno+Dwkigjh0uDEQUQ/9AbNIhiKYfQ9eCb9
sI1ZbChj/pLnFL80V46w3DjqDkJld/i7WsepwsFAvvKAKcXCa+IEipuy+XKTG4rvGBDTUeiiL4Fn
5qeFU3O9rtCc3YAGzsQlwNkw3i8zrBr6wkKcr7rVEbkCtZ8gZx2c4X5jQD4VBuRlMpNhqpuOtmBg
ClFi0q9IYIRLhlG3ndQUFlbtsvvV4KUiFRss2fm1xwcCbE5LYVlrClxUTwOAhgrxNCA4V2JpYVyP
+++5JP65FN/NL63uYqELNwELaJvzR1O8OZbmjkueYTXeIolVqOiZEmE0krcdBAz0r58LLqWwU7v7
rkybFNi7rVao1Km2ci2EppXb5vLrLBmc+iuQUyoNgd+2rRXVZQPakKmL23PTGrYcd5BgOGRykeQC
l77wqh7J/eDQZZgJnbaCQ8+d2FNEGEjWFeHUwiUEXHqZjKjMWnyk5uQ2DuWb7wvFdF/oA8Kbr7CP
0ea/R86GdoX6uahIcNXe38Ja5UBVZUt81BUBAMfdfAc5R8DZ+OOIYYAloH2o/3lT5SD/vE3rkRYZ
vzrP+/UnuCKYn5FzYDcVnwuUMq3PV8RsDWNS1TRFh8HYpvGgtvNGSf3TYLs9knjabeUc+zkMc8t1
FC78kbTHFvweZSF+wVhJLkwzhGSPDp0X+N5kM2nslK0Xguc+uFl4gwEtAqhYyQQoG/Het0+PcmAq
wY1lndH4EXEmhMqZk7s5MUk87HGTuXJupKvD15I5BsnuIBcRSDkdjp4jX0MvNBQosxit5NfLa6IZ
cMI2PFo7FbQGi8ndfWR/0LWtnekY3PCh8hMiZbeCr5uZWjmx+qxsfrvxk45FaelfflJQe5RmEDac
L2rG2qbiMy/bUjHFnrKsrLkea0hjjFVsgGmbSstUYbAfhk3xj0T0kvOk+TAPQ6QgftLWuZp8vP/b
PI61Z0AyVv4q5zehFKjKODOm+g/1lM2P7YO5n50lp1feUFQgb0mHzz7tZaFqi/TPZJP1zDe+Z8N8
0/JbBwIJAD/+oBwLx90uEgbJZYWfD13K4mrHu67XU3Qa9Wrm2Tqnbr0AhaEH+g/ZQex7czeQInAw
3UsDg4Ak/eEK3mPGibSvUTbUxWGQ4Ekl3FhKtNfkGqRl6l1PhbJSc7VBkoLpqCFJIjJ93c4fvIa2
PaKezY6u7akegLRXSrTr2nT4we+q9R+teFsF+ZPC9FFUYcgzWi371wmmEfdSa8bnKP9Rup9GU4It
N3Fwz1KpJQvmUrJAe+Jq05DQ9dhrdociCRpwCrEbxBUIl1Kpo9qh5cy2/1pKtbLBnHwh5lMHsM22
tSb0A5Mtu2zYOfWLQJXPnXboTSF4Il4uSwwkLYiLWZTJVk1wuaLSVy1JVgDjr9xiUwX59LLtaBVD
tvnY7WSgzhXeNKZ/8pNS84rqG/jf4FPhbHTQJ9XXeJfjwnR6xQbOzbQTKknCB2qL9b69ukx8e2H5
7SUPfrfckdR5NWHqAsh8oRVwG7Cpojc0ySd5Tz5aEWHEnQuLbLKU522LEBFzoFagbkpRr4s88pMv
ZsGyRxwE+oT6PWhhi9rvH0ppy7ZHcOkcvYj75d6hdHfmF1ReYGWyoMkvMVXL3KC3LA08fI6tKtJc
fk9XjT49zjihkpd7CNQPGv0WaQsoqOHCiRfrjXu2f0Syt/ccn+fxd3E3tlTG9O6jGa8m1HpHF3/m
t/A2BFkMAHAKiqEXpRR+D3Z8eTBElE06cjKt4B3e7fLsl76TeHqNtCYMGBuS7uo8CTgqjIRPs0aU
086/4/cIYlYHz8doJn0IwnFTooIsmFBxuCKIbTvYFfwmDxvTVNSlOeCd0i9uElkiNIj6zVfOk6YF
b2SBPn7RRSOz0Z/raX72rUZPhd/aWj1uFSqV0Ipsw6bKgrJT3wf2LmiRy6ElMcYKQVV+4SkLicTf
yTKmelH1qZ6qcaWbe6x2AeXNrEe7CYPl9JlQSL0k9MOo+G6eoiELVtiMwy4WevzxA4d7b4xjBGlt
sbhGPUvur3u1dsEF2TyuezI/xmdjd+uX5GqzL+wqx2AcZ+4p2cSxuZIdcT5nNBsU5msAhWQOcMgH
F9WBukJOWXDCnEAtAIDRnmErCwuUX8xzRWnHqvZzSJB4TzF87fqLupGe2R2kWtWbqgpivb6x7cio
nbbfLXRcp1cgcj27hip8k14YHa33a43aSqYoVvqKgxcH2MmmD+ljvSfV0gVe4ihxdHBa9g5uZjVl
QSlgE9I85uVmoe9tJRGy7+wQJ7xHwYiaW9rer9CdDJ4vuO45R5nqZnTJ6vt8zN/4nCNiq2VzwNmT
UOvGiLljk3IsT9pWoEoYANw5npTb/kwBCUk+zoAFThq9zcOHTy6wQ7SsiZt3A86CADsyLwa3K2fA
BEj42w0qPbxdO3dnoAkLIpaF8/e54FguhQ85ev3+i99xb/FZrDMDhMLncD/By1HrtuHjDr/abetp
2JXrSlzgQPZzjfWOgzCPO3bb8FTooD+CvjWDOUKZCC28A8IMvfcIcKVv3og9g/7iprpAulOQcqqs
edRXpZFu0iEkuGZfsylf6aL8/N3Iw3uoSL7iDB208R+cNc1P0ifHKdh81OfLHkAUjFCPp0gxsEMq
WrBRhS2IBVCtP0rJ2sQSDO1amyZV9JLHbxLED/PPanomrC1AXcBAFcGJV6W+HkIx1YD6BKRr46+C
8EgicTd+nA6Ezh7Dx0O91LR0gnbdWH1Xre3NY8CTxlz8vH1GG8iUB2PBtHsaGeOM7kFJxWG9roBi
CegmAluMGCT08hlbHh6z2jd8hTffJ9Ua0FrQ0uYjehDTrVvzvM8L93Up0LVFaN8dq8rBX48NUckv
UNIKqdRdj05lO82XnLnxTpermOQWqxW94KOZfNq9S0uFYsmStBeaNk1rHaMjh0v90/OiaMt1XVNZ
O9gQ0f5XCTL2/rkhaWKGOEZxwU0dFREcHUpxckocoJj3vtiqNO+Ewr7YWIPEpvRSldQtUzFIppjN
JzvrOq6Qy+xwdJTt3T4FitmGpyHoy4H/LYAvZ98wmKnX+TYreee69n2gqES4K/9va5oACyO1lZUA
Of9jkuxsExTgCmeBs7WU+SLpo/FYVR5IqQk5ZrYG6jcZYqy8blP25H/zqHObVL5aOn0Olj5aShZs
bqGGEiPi9JhN0dMCz3IGs9wRUgLtQ2o/TdUYic2++FLm8/LRlCSaIdT0DrBG/L5dLnFobVT17Lv4
fu2jfuna1HG2+7xBvlBoPG8NlRVH6gDApwkTCnavm766vC+kLNkAXCeo4uQMFJYy3SCdgfOYfo22
bIiOFKa36i8F1Xcp/wpmGOQRllGn+DuBVwPWe/rM/WiVhkNdlIUQO38Hoyp1oMmOMszYWbiQSeQz
u0/5EcVVGvNBRgAu5AHGIIwxuoHFeohts/twCpLZeOR0k1F/4ZMRtuCYF+KX1iVK2+9Voc+JCExL
E/PVqXG1P6reoPedou9dlyr1jjaFXDTr0lErT6ff3W+8F3kkeRvKBP6hnX8TnF/D0MzhO2qTIpO1
/UsKktJ30RIut2CxmiZtF7B19gR0fYlfaMJbFZdytM4uhH2kPAoQXXGgFjk3R0dTrcph28HTwlLC
5BdQUHXPP908NMcRnZjThCmaJkTMA22HoGo87hdv87ef4SocCof/xOVInQM7gW8SMNsA709XUgjZ
K8EhtTH5qekfUphtfaZK25fVDbaElSE+fLvYskWHBflJcj8d1TnuuO29z4sUKBUdKHknXUGCji9h
kDZnv6bI7xkOgKO9xFazB2I99omsWdC7dB7fvMU/JSNBP9dj+VdFjtv+iUb+iLeCcPaSMZKPJqd2
MzxGzjDaB/zQkzG2jfmBkmlkpEDAyj8MuwVKlnbg9j7HSzRGZ+XDR2Z2rlGn04E12/0OgfXrLLKy
qVT8NwsnwQoi6R9XX9hGXq27ygw3BlCFjbXd3ZRxTYG4q/NRc7zD0OcVulp+Xw/dS16ljSObuBOs
y0Vf1BIDQQqUoGlZViNzj+4wKfzxS/n8yhUalb32Ic8jduvSGboWC+GDOsbP1jaTcE/g6j7Yxg50
VZWzAT9kaF5meM4AD0ixxUfL4UAZuQEeQEV6gdCdQDkj1VlS2FZKOOIEPWK0jOfB4cIEXg96/5am
vpy5A7ihK7/CltxfJ34PNaPRzH1Qo0+tP5TdalJg2Wt0KJLP25IA2VB1itZQocMSs8niLiLq9TOq
k1Vdz7RTF6BkDv/4SIvEaV3P5Q+ie68EiIyeKc5wIlQsj80fDB+LfNepAdUXXuA1R2bdOtyKrNxj
eDoZkqxqyLCNy4kABPJJe9zqzaz9u4bkIoXGPIIjt/YnI18TfMQW9M4uEk+mQA6xo0c4k4oOPXhU
9D9y09A2vuXfHqhO4Z0sej47LRJBW9TRAnc/JQGek6t1UpNj5T12T4jwEa9QI0LDNMgAxiYceJKm
jXiY5r0UGQ6tc6OBOqa+n0T+1kj2jQrozaWQ2eFrPedggFUqIPThVYdFDOxHxiAyvNdx5M3bTxk6
FXUiex3dzT9id9sgrFl/RQQOLLW7sxyzuaEviTSsbJFCGNz29BBttJ4xW/T56vlmR+AdneZc7CMT
x02S9Ln+a+m98K2uIrxIBl0y/zLeVEzrTVa764Zzb2eN3x2/P9pSD/GiA1+A6yPaO+RwDDFDt+rm
XYFHczQtZ/4OsG8uk5b+Q/NRGxNPEubx1BAIoGNEFvjIqs+vOJJso6Y4gqGuve3VBfJ4JcykEpNV
dUdmz29inmqBlQlajgJmKrUdE35ARsIKytyS6jyX3LZJE9jTTXSmmh+FtSDx4W4yVhtecJeEz4LA
TqS4IZCN2xNhEsd3LrCxzv31xP0Wv5IQNDTKFGIwDRxGi4kdwUJvEBhVA9GGJ1e2lydKdGCF2ewr
tg/2+qAPp77pbrEKlzd1vqlD/3bdRv8NzyReyy4hMXx28nJFPhTXvBzu1v6IzPJ7s0tLVtPp9Bkf
zO2UeoUHmk7FCCdDKeQne09uBZeLoZNg2O0mG1lGvgLZEPkdp8OXG08eqfQVn8yiVxQvfB06Ges2
7seSuqdLGtvDfGq60LVUJA/QhXMMi8zhOZOmiWVEz2hhaNnsYkolEGVzyw8vEK29k/+C/fn7DblO
1OmBCWSdx1ZCLcoYAo4sMCpJFXU3IHxnbWQ3ZfevOz6YF5Gv6DZOr4RFwNMYXkg2aa4bpoVtf4EJ
EVnXmBQ0LoAuGdq7wL9xW+EZyMUBkcV/fmYqI2bsmG12WDsTVULsApNu2OVZwqmE47DVeGDXeVJP
mW+Aff2s2Ialwwqs6lIebVlsNC2AxX+gkF3w8SmgAxv8ydl24kZV0UefzTyHFFsUiMzlwX9cyQMQ
q9bLVJS06xtsu8uy3KEIflX4l0HO8ch1b/U0sBl0VPEd/5+T/kiC93KGc7kvrbmnT4MzZZBG3ZjX
A89OnXHybVvTLZgd/lbF3yy9Fkhr4dst6/y68jRTNy2Ihof1ldYzidyI/JXD3tup1O6tJuAl+WN4
scBvdD/0JEdmdwrrBUkmAq47iS0nG3CwGLTZchuWeJRGtwQOtFMgV+w5FI+01oiqm5qzm3l0rpiy
YVqTGmu/j4/Myku2U8vMB9jYjhxE3SdCZcPocNGiJMQk9B2pGAMzaKNmHDBPvwCBAe0KENP9YvKr
8v40Y+YiN5xwZ/eJ66tehZgDwejxwI9g2BfGH/Au+WUxKr2ZPiPm+xP7+hyBF+qshkkiqvCp9Btz
EOSOxU4HXPACeF3NYcTP6a0SfBgwchbdXlESDC61jNk8jg0WTCp2UIJPbQ4wR0jpkXiFi6sWZ5wC
bDjqkwFGG5pippas8ymvktVmNobVP/yIZljS0zxeBst7a54HdY4lNVoLLbrhTVBzLTXvajEq6sYi
jae+E3LmeOPQZ6f3UVG55dkTTyxbh3BFjReaphK//8YfrO3bMJntgmLdBnmzmiQzU+prYGPIGhdC
TLRGi4L94zNxGdJnw5hA5A/zPyume90ZC4gJHFccAMS216SIF2pjzwvRQ08F5JtnmdX50YlLvFUC
7/V8IZrJUb14moZoIxmWuwlvkhBQ/ujLRQpj1jtVEaG4ONFavn+lzoDGlhUeRvp7EtZD7tsoYBSy
rixfDcG/hiDai/Ri7h0HnY8PYrdSFxAvHEhZ1xFaIKgeeoTQAzNgdkZ34JUUcGXsA4S/HKz/FC+H
MKvxnl1ZREJmz+qXyUEZL5uibX4iOlz1NZQ3671eUOldv72DjXQFqDLsiMFNoSpTgmp7Ob8dQjjf
4ww0idl+eQLjHVc0UJBpteUc6wIb/1r6ZOZGQ03n6Tvcaa8XQOuJH+pf+k4nsK0mBIm9HRxT93nZ
9NTv5BDTQbqvlTjCrBwfJhwd/BFMPSFVnkEsk07ITRuLHAeMpJSYKti+WA5zGjF4RbvyFaSLYi7W
iFHpZx/tU3OwuY9XyfrBrOjcSe0B/HhUQtVbhrs04CKD0e5aaeR6RAticSgWQykwqZ2e759bAjWf
qr4i9Ea/5UsjYdg4xI4Gaazj65nK1whiBzcTNPJPH04nkKln4KFNFbVib6xZDHyEbSkaRKjnTjxl
YChC3toYUio3GFF970BodCnS3Yek5PXOK0gSnUawusZiZWZd9GEqJUd1F8pne5KsTMK6w8d1/9lh
QhXwDS5yw2uhqrAEnq3civOImxohf9J5XGS60GmU+X7jJ+T/BZt38MDKW5IxDBRC7v3oMhhgM4gQ
q5x+0eK9kgeFz9IL0kHKZpuOSnzO2SRsVehi4fR6fzR6iNhGrvS592s3ytx0KHZhOYuf5/RoLrvv
X25nZ0cCQnTOcmIpAgNBt9aw1xNlKlxrPVAM20VPoLJei/5+F75SZFEQHMDe+0rzTcWSFjZXt3EL
DKNNf7pMvwaBl5JR02RTG5shV7k86FkSjQZSyTwpfw/M7Yz2fuOzTyMg+zK1WKZsHOwH29MsNDFt
UnNX+QK+tpaJFGN7pIngRyArmjyOZ7f6JBHhFgM0iWYUfH8MJjIx/rYvh7zT3b7ppZhK6ZzHZAaM
V//q8twkY/IewmffdIGa1jCqqw6HQ0GrrswHvYXRV+VPGl5XVCdjPsrYbWRTtjlh7woA/Ar46Wbm
w159CKgm3kOO2ImiuDOuEPXwRnS3lSkKFHLjUBcI+jD6tTXoZYGdjqaJySSUNfzvmO+VfRJpKnOs
F2xJcuD0l17/TOhy+skA/CSrh5izeYLB+sPqx90GHElC6mb60c1GQdvLVBITLmGrhifXTMqsdrA0
hHUxqoJzie0FjXU6sYCOLKYwJARTaQucuT5HAQ1VIBFH6Q1ATDPfwHyNtxsvzKCGKYb94LJOGoCY
ZX0PYmXMxyzlZQ0K3N0GPIZ/VEsXHcQSLN1Lm2mNrvVYBC4u3bjj5zQeyqXFCr5FHbZF1D/fF45U
MFmrMpcVJrRgevGvkR4F9hBdlV3M0e3GIAX7Ku2RuQZWBEpiQb8B1ExiEOt5Cm1YEaHJ830UOqUa
LkgSMyYsN/Op9nH2KZcNYyXya9NL4MkqELSr301K0UlC6QBMK8o5wuAB0aYf1GvReM9MYLJNOccM
U9npmb9X84RASXszyghrcKMc86pf+iWrLN3CqU5/kWWeAC09wS+CH19Snv3ruVGQMJ6TPsmpgaMp
mj4yt4kOF6il6Zfi6JyDn3dQaYAt9HL7/FZiDoiKrd6NmuaplZYJ0FLreufzU3mB8PUJoBS1orpc
evlDXCFTcLC0FrAvWjXbuVLZn4lBVFOllP4jXfrQB9JmDuRoprk7gzjnfruhRytK/vtf4AFxHMTF
lV0WlUYy7kuyIa8L6NaGZ0U3EQtGeMqnmvcq2xgQsr3z4o/rI/TrtyDX8DLL3resmvHBt8kqFWYg
NRGh5cs8/h79gJ++ZB3gOcWAVs3qRN16p+I7zeslrui+VWrtPYvLmSssOMQOMeWDEe+zx4pgL5lB
btzPBg8oGog+9C0PB6R1/7LPJ+qTchovTZcTCWFCsoaKVHkvrqAJuIuU+Y2Nj43TbLs94Os+J1uY
nvqyg2bflIiITFnUJNOijWlqv2pnWMTB+EywtvEPu2gM3vlVCcA17UiEF/3+4pvRQD2ly+N90lh9
fdNfE2Kldgw2nrLQHiKtbfQ3NoQPYn0MzTnQKpjVAY4S5FDBCqCOeYmP5mtV9+6gAqivSN7KGc1r
p/+aWfTNgAFjbEkmMyWH5eClteMy9jH+PyioqWpvIpp+Ew8WPedhcxaZFkbMsYClmjkGI/J1MIwL
tHnmg6DEK+/A1WKfx0tGGM8ymfY+bXLyoKYFzAeCHsJrDI2YxHLegcu+pBpSmhRJvgPcVdYX2AHC
HnTcbxcdjSy3caMC1iqi4ib/gcRB30s53c/ksE+PSrRIFEhm17rx30OiO/J57p6EHVvMe8caMI0h
uJa0qOr2Etnrl3wSzaFUHmypayT5LA/lu0Hy4d2IMXr0GAgJwZ/U+H4U6jV0w2UBjhfqsh1RxsoO
lPTiFwOV1m9WEKuJPnF5g1RcPgudLBNTJ96jRhh6v98plO8Es9odkLimbh+7Wnyx1fk3y2Suwvg9
he7TCsE++e+wZrYtNF32234Edq3gZlBVeaSVxD8Rw5Gl+35EDYZBcq3m+2Toen+H96fK05S1o3D6
nmHJZg6gObHyZFAJ6Ub72NyUICKoEHVN4dI77vp58A9dVJbkSGMgnCVTBHnjZYfsh4YmYCa520uO
RFcKYVCS8rneKevdx2AwSAojsYe5fMY3Ib1zJqc75sB6gR9HE8en8n+udVOtS6pzqnoissvjwjpS
ZEpmTncRDWhV9ITi60Sxpk697Op+VePy11en3UfZMIbEU1ZQ/U5KoEBeuGF2PuqIj5EGSLoMR5jn
xYwivRWuEpIToHCRpk5qHK2gQPsftbpDin5P+q3E7ZMg/iLeNCVGIBXcAut3oU0iL/cVeENT2nPB
yKn/aWGjQTFaGIjFXoMzuyukJkiK9kJTvGpOFB0s4ey4J+rtWEceeqV6Ccd7RUl201U85aNE8mds
XnLygRrFHa8700Z7G2HJrq5UsAfO2/B5ehTbVot22GOVBsdR4M0HpCrG47TEP+VXFID91NPVJ2Tj
wsWP6XDgBXTr7s/0RI26XcZJERoOo23H6IifWiZbgi0MLvVKCmgnuOWRsIMCGRzerln6Q4cLy305
evGI9zOhl8tof15oRfVkRvkYAPmFuFRd1AONzngHQGufbLwB3bLs5Io3l9FPO7SkhbwSanxMxmqQ
6JkbsaHY9M+ltve+vg4X2Nf7lf8U4R2F5h3nBnUUEIBvzt3rQH+Wuv+fn2mQ1/n/zrD405Df+Y6c
7h055zQKUUsOghdqwoBgdNJSk3igBZsz25S8xEP5cx5QJc7CmBjz9GOLqZkCMU5Eq1utvibPFBpB
zME68xoi4guvHzirSu/uUqUYp8yrAxAJiU4x+px9rZ2qN7CtwESCNpF4D0NFQmx3RecP1eRR4Ybh
ZAmOWCDtjN6wnrxTcFLV8SSCPnw2vjOHaC1m6hdgeXUCnd5GUFTuZmziehV7eJMYuMrE6DMIxsPc
CYlA2KXrU+ZBnSaG0JOdxnAu+KJLFIpL8NtQkiU2StG4UqUlMp5SpqpmJIIoNshl+QQauP7eBWBU
XlfU20+eAXHl4DURx4tQvC6I39NAP5SZdD6ehr2iDKUe94g3oAJFTAIYbcpwPDzUxlUbq4znMBBX
NAAE+sGD1PpZFeDLbZ27vm4OFQI3NxAoN9C58Ud7bnxaDgPcBnj21kovkVaggQ4d2ruZ7YOfzNUI
sDLtUhdxNDHYTFM+7CXBTpBk5NYM5OteeRw9CHdVmnfDVs7AvUiBC9uGhkfc+wjqlk/UXqf21yTD
sI3yC/4xl29qztFGslEZgsIucDqJsSD2O2bG9OqqGHl4hAfnkEp4pQU/wvqYkJw9HToQfY02hHeA
sn4sQwnQjJPkovwA02pfHn+Ann6/1S23WDdIcN6s4D0uDvQCArFloxqrOMpuX82uJtVNL7kgdXin
HnOJf0S0l4AXBUAbsFCewmpU1nFkjRt0pE/VXAuTSiy+PrEV+uxbjwOC2rVuTfdQGCmlUOFIGjXx
ftRIiWWVyXFid/sP+rqsYEUuO1cTuwJohJd/1hWW3L700//H0L5wSNLqXjNIIwR2AXTMoM51AEdX
OqiSAnu/kh6sQ48R1dCVElmlKDuAdhvYtymhndt5ruWa7KtEr6zulg5gpVKDYRKOXPumu/ATJTbi
Pbmn/5sww78kLtGTYak+NKm6K6vAFwLKvqq6Zn6c1YWqHET3MNCeDhQWzgtP3JJ/baYxmkqXBOlf
oXLiESDcctrCmoX0zAnS7FFNMA7DDEvI+CpjnjZh4qmUbZlYsrTjAdLtYivyP7anA0ETKIM9eqCZ
9yno9J+q46ztPF6ATxKVrOnqjm9wpZuo/ZtgJy9RWiyWA4CJTYZTX+JIyL2AJDN8WGjasOD3SI47
nCD/yiO907IQqViYDcKWSqJGxog0QBxIU/GSRaHt0/BlxWs1A+D/Ybxgxwn3O1e0tSfKjxZmzgF5
9hq+PL3SO1nEjiS1/1dprYKgeuirEtFKEeGPATYUXtn8hjWMEoPuaUbQXFsmy+fDdcYzXB9iwX+Q
e0d+CGdC6EGRy/FYSXJCwOU2FHdty7CxxXVje5mXEllAWerZ+E9/KoBC8vtKhfg7wFtU+FRBRvK4
cWSM+gH7ZQawMa7ALG4+E5RkJGDv3sAVOoCCJwDIf721e2l4LlLYz6zwAUkF/vdnmXtk3iz8zOjy
6bMJItGOmHEKDEkDs+AxV3GGoCwvw9Z7h8V4zimZx+3CpiyJaQ8j97M6m9HpbW20pYOYCcnCnWfQ
m4PvYZVwUhQk4XUQ/zkrV4KbqsKbVeM2/6DElzZLQuX8JTfxM3amj/7UtYDFbJ7j/9bNrq5AvH7J
/mEsNe6QgeDgBeYoK8QIKhepRXSlml5SopQwJFjFBumfL41um8VvJhOt/NerSeLJCLkW6xV8ys71
JgD/QKRhmgT6QUgM+vRfu/V9A7qJw5BMgCchQVQMF86c1ZkOQOXJ7LcsivckYsorUtQHR7w7Xqxx
CwNLe8k8+izvQSK762v+6GLnZWnU/p33VGjH/yps8rllVBlL7W2HQd6P2mQcpgH7NnI7cQsYx6dI
slxeA1+pvaMk0hK1+5KZjSybfRtxt1jHT9nWi+7RGB5iy5VZX3x6qaaMPqNyDPzXh0pN7MDonmLi
IET0guM0ak5xQo5KzGniA3Ob4vH9ols2MCj7r8tgt5M6pceGcNeam64emCLS0ma1hV9Bw08ZGF5b
5PtHYDEJpu8mV2SllWuMbWqGdMYhoD3gYH4rE/kvPJMHWTGtM+NA2CL6psiMQQ8bM5kVNlKF2Fgx
lQNASbLeKJQp1ooeocjTcA8alEy3526rDwdRu2S85GVVoKsg230Ewe2oefNFXE/yKdEWvwS+yuWB
HSxpDSN7PqMmaqBYKSWeiIfdfALDi5GIfSBSAniu1+Rib90QDo2l63rZBr75dlJiFLTkkLnyHvfd
D6zVI/D5beaVcQF/Z89vz7P5HpRtJuH+JLveiMsIXh6u+5MGq7yLXznlfO2i170bEUxsBp/J0GkX
aAUkozhQ9Tj16osgzfrPmcAunBkiLmmpwXCOcMA/Y9Nns4Qdsba/VVDYhuXEDb10CrquOsUwobFC
ekr18an+9kt18QAnlDmiCbqWSEDOMY+jBvn9NthiifaphEyWC4rIqKT6tuylND35vHZmfhvXhzOi
Ndb4NSk8otNKYLePK2/8rfMw4WzdMgwYiV49J0ycpGLgpQPFx8kbN00eE54FTzxxwmc4JP7IO8w2
YQn7PR9sX7/iunc4RyDok1NDYCO4hA1nmK7x10tU+e9zW+LtTKRq/S+gKTbTuo9tuIljAw/iPmrO
35M3AuJjPLRiPCXaU9Dbl0bcmx345KNHGXPS6tj/q5BqyyyndcIQPIhNcvkqW8BddfHgmbJIEWnr
g/exuiW35ZSl8+6wJJovTylp6vyHFun1lna8Tpt045JA2bMuELCLHJ0ia5Xsndyw+DiFKqeniqgE
i9Vy71/s+3cBXOSXiP5lP9P03dhgIFktHKJS+afMdVAfoWNGHtQ+iIQDMKVzEBVa7v3tyteiadwo
nQG/1hKz4qna7dqBIZutuelRyAkQKkurtcPJOgTPllr6FnAdZ5BA5ObQPyr/GUfnj8Q6BJ3g2RYO
hNjUyEJliMLPaMIbDG85/oQkveUrNfh2Q5qCQQMLoyGDaLY677c9X4u7S5apzp8jD4USFVb97ulR
4nxvb6bDB+ayHAVkGjfvUpNeDo0XJl0MhyE3I13mezBky/zicXy+iWUwuoUy5G6A8A6gV21MvF58
tmi10915RS/3ffmklmS7iccoDoGWXyh41zBbNne+FBfSV9MU5vc8RsIeUecJSfGSeDhM4KdJFRKT
YGJD1DCFKUfLN9kiQl7GVFHk3aXgVIC4llhdpAKyGyrMFZfAlV2tmJew3PKIvRwgdVsryNrtyPsg
lsy7oOscVxU0ezlt/Kv/a/Hf/Pj1S28gx0EoITz5xO506CQ6vCFlfPdl6CoY6KByPDzbvc2DI4HO
p9PmlAWGqbazUABZwqEG+3Lk/nnD/zE1GY1cIM8CNAmPfCH9t+dF0BpynTOwAv3tEYQ26OjiYyVZ
cBo1mYBpIuoUj/p1pnoU3U0bW+cSWoMXp3e7Xw7yjZCUhricO2uKMBR4TYMGZrqgtW4MwSxerwd/
IcAfwoA2aRv05tAxSNsjzvfFIXkS7Munp7Fngjg8I/arZ8xo3nd4Qk+pyMYvxeXN5EF513BwdMVU
jRWCVVEZfcNUNARopvdkJhwWAiFczFp10pXBmErJ73+4DSUF/y+S5qnuamn6WJxkdFFF8TetlYFJ
ZNt3B5TeeO04tuS/ZQhLFnClINETPX9jYQ+daQxn22B3tmhmRCUAxEgTCUddMqXBGQuS2WW5m8j2
ShrsMDTyRGUCqrHna0SfMz++tj12X2V/trIwWjuxBBhGZsFVwasyGXHd+fhYtXJnzfP37TexhxPX
hSZn91cq89XyvQDZ0pFOZ0mbWwyyH6Ts6hyR8OAP+h194f8QvASg52BWg3s4Ci5MGE6UiaOD1WB6
Z67CrvlnuRT8laUaIibyZykXoYtukpqk9mUdDsSHBC/mdExnMYQhjIP8D7TO8/md6aAEyD8eLJTO
WkjY+iijbKPG3wwBvCzpsBc+NW1Y5SLE8RRCrx9BNtItSO4W1Z3Qarq10dV5oMvMecLR8MWFFOe0
ApCk3HeD1WGrZM8qOaFBcGPAgMV63ribZmNvfkH1wVlpirmjFIdGddzQVxKOC8EKqHHnBoDXV70N
8ZjHP3Vb+MpfVm48MYjmMYejSe+wMznUPjeAbK1hkjeJFqnFbQDi2f/GUiz/aZTWfF/oFry1vBK4
I2DS57I8LYY+e+2dy1JMkLt12m15if0iiy7apUBuPcqxYsmax1/Pd6FtpTpdwbIB1T0bdavCkpua
Cz1yESWWju7CHs5VDu47QeoelToFoOCmEeb2+ztweh+td7T4aLNYdAhiEscSaCkXsF1io2xdNMKx
K0dliaxsvn99DDcmwRe/n9GbFihcAbJEGiexx2DD+ZhI6oanz647RfZafBFz20ALE8BGJoIk4qul
o1+nWyBj5NNbbp1Ud/r6f10PbAVHCsrYPnMOJCnuJT5X+NpP1uxAZdGhRTx0LTE+eK4ghayji9lH
MV6ZCl9MMvgAWjOL3OZZsOszD8zF+YlEJdw3HIMHZx/GWWSqSsZkQZ7NT0x7PTkW7pZctjmj8QF4
wdyX6nplgLfO4dxOHL7XPncG+mQRZRD32099//QPt9Mv1u0v8Nj/dwkuyzaFPizHHprm7zOlKdPl
Ejubh9n8sdoQ2u/EzatmQiqo1RD6zp5xz4BEmpxKx4N+5eutrYiCE+zrLm7PTUbLQ4OysEvC4vZZ
/ZsoAvg+AJSW4BYiF4bPz+CzndzjjeN+LU9wdW8eU9S38S0rvLAJ8UcaAj+fPQ/pNtKw3L7vmcXt
IYQiB9ZDgZ1Dll7NI/jrgGiEeA6h3qc7TPrKlLG9PRkpz5m1/A4OPZ7NPoOFozyIg7QGLwBsMxh+
XEvQxcNJE5i1YeF+rvgKCUm7LEnKkN7oFYpe1FUYlp+VYuZKr7sp5QE0e2Fm+3Yz6h9Evjoc91tk
nbKlTRlL1xVsUYTnDZgXmQmIq8eZDi9bYloMu5TTx/XsVVgL8HoUiSG1BFcET5uWXiqL+NoyPsKa
DfbWpUNlPEiEppZ2X9FBNgVhbzAithuG0hXz1QeqpOWPRQQWqvaCuqZCyf304Y5/JeEOVvFjiS+V
Nu6Wsz/CTC9gQ+JDnR3BkqwxON1ZKExGliYoYQVUvitJNmpdvA4mxRENa6r2nlYjtqkkFVqzKSIt
YqO4IDtZksZO722z+x+xIN/+UT7mcob44uCaMvU10cWwfSMv1PiFMWq9ND7y38Zxu38IcTAvK0FS
4SEVsfvRexjpDkB2rvKaIYSoShpHF0b/CtJIOBGvwnRZO2N1D569/96vcIncyLdpxRgB2QQFRoqR
IkNnCk8OqgL1tIxZWEkur74eVdnNwBaTxa9QGVvg5aQFlDLLhp7p6zEDeC+AZwxauJ6p5E+HLUnz
feAhp/MVjiwOed45wHnN9wOYpLX6FYNRG15ysKCueIzzsBPXga52OUgNBVjDvzhNkJmtOaE2xqqd
iyoF8/sNc6AMzpHXKA966dll+rWtMcrV41hDPVkkVe8K/p7R22ZvuG4+6KiwP6qXP41z3bIiP8sk
KfODQ40++EZnLMo46DVHGIBehg8utx5isuALovUzW8/0D7mI+OAKUkz/aNVfpQWK0K00BFQkhDt1
UPg2zTEWD0ZbPxPim/u5DBWya2CnZOjcXuj7weTPEdy5wsQU/1Ae6JwTZZcLJE6h4F3lgPNnPsfc
bZf6uRFFUgml9ZG4RX2Jibk2v7OsYQHqbvt9+JjouUt2cKuYZvVwVxTvYoin0EunKZCLfbaLrl3h
epub6KAJC8NxY8zqdn6VgTbVmubVn87d7GHN+sdAPjUzzbISfv/Q8+rQL+vfeQ2sSXzn5KiLnsAX
MbJcKz8o4EHAr6mPlLaqkLsdcvOsh9xMmLXNjTi6waKPp5G17aE/K/7ybcBiK9hopC7cpyad5hdg
rkjwqgofudO+lMQEiyRTyTQt80JjykRhN2vyPs3tyoqLQep33mhOII9qefNq77UAoMkf+RUeCe8m
ts2neEUbZjTpJjpQCqmvPTMRm09WWT8+pBP/enZ7+MpueburE4zd7z72EJfAw7hrr/ZdPMVs46OC
JirEzFxYQUpka9r4RAtcDHya74Ye/HsPJ7lCV4WeXtUNMm/AdiPsTaPL9aGC8Ylm7nG/w5AcQQxG
btPJ91J7ewSw/e+ZFxJc5EYJJZrCURBFWPvvjV+HalsdTvRR36ou1gkYujSDDPP1NpAQ2iaK+rgr
ojkWcczBCB+Ew5V65z2oTHud97QgZSUk/gyakboKUgX5gSMKn07FydDUJYEYBEorFqW/Lq9fOJbw
QbG8ev2wu3zTzsjX3/XVYwXbxNO4LFbK6qtU6EAPwnL1zBtlicA5QeqMpyrOeC1MzLveSXyPeKnr
hYa+E1FQbMDbSaO1+6qhbPR/fl4PpwkLWW8okBg3OH1uM+v3641gyTbNSzGlJJMDWT7BG8KAnuXs
xe9RLVVkRIMvq80TgVUE2o/12XRUgghOcqa8ZnkHpLaMvjfDVTcamcuv23NbIHL2m3yo+AzT4p9p
Cg3HBZQ/WSJAzqIiHb7yOwKZsLLpI5TFLlk3UFS4g9XSAr2e+rhpSEK2xqRjhmV+U7pf3BgJnipk
dhquatrxiS5Hnw6ZOFyvYWO1oJypbGAYPpCEvHRAmAFlOypruiG/LKaH717ftUM8PBsOUDYOZ4dp
QLnJwxw6jvPC8gExqFeK03UESE6eQQN+ZPMwlYyUyIVEHcNIS2wnYTBoT6tVbu2btamvg+aTPUAP
lAt7JVJM55KxbUVr1T7PZewPb7+iSDlSz6LzlzIqOlra7x2DB503WAmUN7CSzBD0kl2KdaVTEfiZ
0xJNg7L8+mBju11KxzSwg8C11Ks1fh9+iQt47dXOt44IDRxUu8Y0CR5CzDeFmz1vlIrQ+TOPUpJO
CSwP4LsPilSACch58rSrLU5U6/PHqMFoavjF7o1IqisPSP46YU/1UqdHxh2z5kbLGw+XhNkL/V26
JIUZvgRzbgKo8rqNhaj5Oa8ZPKQ7EFPePTImllY1OnGHw/fP8J0kJZjb7DI9izyiy+WW6lGABtt6
fzhxsFZENHjIExwTYVTnz8RFvlQcoe6e//fyGmPVQDURHBqHh9xYpJOwXc7Cn+zTkBUOKaAOrDhr
DCt1DVMfkNEgOFqW0p2fm63CiGDwqu0/mzDoU/jojjHWMQP/8ZYw07JcNPe2wcmgodE0VsKHb/dl
fBwjxd+KggMa9HYi4X/HEew3S/mAIO+w4mE1m5BV4dpRls75wopM70RnVDXC9uMnqGBAERCHVwr9
ORPqWlWFZ5Qt75lU4/L6886zo2Ml8uxM1ivHCcJs1BoRQ8KubBASDsNwt1m0sysKBXWc8mxeCfz3
QCz0shc/p6fJM+wbZlAKDReTJ22+ivfEsWNstdf2tZ3V/BHI2N0ob8h91nhntjfo5qoGZrCTn7Jp
dl0saLpgfKUMIzh/ZpW1mUTVG2cARN92NPhZccuT8nG43dVbYQzYPeHvCMND/pgN749a9jLfY7RS
eng/l7ti8IL37BSEpQBj3LMJ/CFojWxcuB/6d8xcGkTKKoZgm8yuUa1/uFcAO6enp9Y2DS1c0H/v
hK8fWzpcsis+4JPrArLT6hU94DbLV/18HRNeHaIJiiH/1Eer0bfYj33gGzynysHkQrtwqFuXRCdX
UVUCwp8Y9+TzcSt9qVvsecEaDTUn8w4ZN3VYd/jZN/PW/SRzyNXIgHyhAeeYGtdM/jA/XTgUMQyO
Vwvhx8KgZQA9j16Ca6wqvtZZiDx0wex6kzIYa3I1tc05biif8Ch1DEm9sKaBXs/D2KBIaA8Tn7OA
tNO4Ldl/tyUUUbMK4XAitYyNVK8gPVnUUZZirmpsfZSOJlHSPPrYhugVMeJIXMcPcNwymZXVcu42
wfBSVijptHwGyTVSOnd4h3pu3z9gu6zRdIS2qvcPPiENWTRgPYr6onqlOtzQJ55TFhgMP2+gcN0O
RdW/IMH+j7Uy7VYQVTvjo4WYfzMfY9r/rLD8NU/b/JOxvQ2m6x4dzobbh/2mTICFQc43yE9Fl8GV
A9+a8qURwnqSxZo6H4Ca3HuPi9F3CDy6KvqemIqCQoIE959PCpgADKA5P4vKzKIn3Eh/k9B+dkxi
gkfDL4eWsXN2SZn39zAuD8jSjGJZvPYQMS+bqH2VAxeMrtuK71hUOguqQrlItrGBS3UQSJsLF8i+
ax86QHEgPKLAbf9jrwQdYZdVzmq8K9mN+maDLCVGcJ5xw4r0ku/JGSjW8sc6xj79hPZRnEzgI+MZ
BAbChsvI1XqzClWaGgylYZY9S5sa7fYAuxzbh4kThmTZrMAECWfby46d2E7Vm5YcFkCP7LPPDoUy
9PPAJO2RIbTALDiiHuL38CkUNfHfFF8fzlPXPd8T88ZKz3x5ZSbmiKKblD7ipteHULUEYR7NEaqW
1j+ZqnDJmMzkDRZpmp65GtHttwdBjI24vOmFEJZprblYQEQCfiesmBGkBtfOK8+iE7oPPLf7Vlnm
SHzOVyOY2PLSmv2lproF+qfqSAnUnaeC+3fT69fHUFj/zXJJ0h5NNsQX1GWdZFT1L3/dtHO5M6ar
/jdFHCPXyikXagxRfvGrWD4dx+ndx6MTI+Ej2HDkyAlNMib42UDAJ+xfEhpHV0ByxKSitvJE7iDQ
E/SHwqlVvAlpqimtv45aOuoy+amnnINc+zyxbPGioD1Wm32QNMEsQWTSkkdEanHMYUz4mRQ176Ia
kMtcrlMCeIZ1TQJyLn62xS1+9BGLsve/LDsAo9u/aAoJyBjKpwS3EEsMqwbDUM7MNHWx7bvCU3tZ
9IQ5g3gbI/2Gz6hbwX/7vWddY8wkbP43gKAuhJmNIWVw2KTaPWKxwRuRCun2WPzh9En0VhXGp/Ob
By4XH9IrZsnPdso953NenGngKN8FqmnuGHj8Npc69LOuEM5A2G79GxWmtM0bX3TV2mAw10WL3RpU
7jf/C4Ob23yELKtl2BvEsIU/2XIplyUHKRYsYCsyzmfNLL/CfmEQRXEyHOhAQZoBmtavb0RBI6hS
7myJnUx9m8zarXveeF4GFbqXgPGcTcBuebxL9JgjgqJGYTY8mP2zisG5PQ719lXPHul+WRbvmDzU
06pBpiiCj55x0oEDiOi6awsoYxMDnLkZ/UeG5rjGbgEp0OQOu3nUfqgVNJx3td4vpj/86FrC83EG
PNQmzZ+JyqirkCXIf2hVsaozoJ+xGBn3eUbYRY8G+EvYtv3tl4wilH2gibsRSo68OLZLuU/0DnKm
K6aKmThzoQYQ9HN4pZkPsb2pjg/xQUF5CZBsee7qx5PlJVgGocsUR38ZXoCsagRPT2s1FK7xpBjx
bSx7sLqf6LLp1cRlot/CANw68fYZyBR6bQuKGWqqca3caC/6oGxHjLzowiUthbJgLu0b1Rme38QL
L6DKzrtSJK29lCiy9lOUdV/IJYAfTZc6zBBuB2j2gAtb0YCfx/wiNQyzHAHTyMQfd7T2C13GkfNH
fJXxIAPK79iVByAVJqB/UlUicoj7LEP/eRBerYnAB/rIpUyXSIZUemFhhj4/6uz8+11ly8UqxoH6
BLMVm2faSGCzIK1PJajk9OUK6p1L3DV5iKf5snP/wUtUVE6t+/HG+Q1MiHlbgAdRQEzSdgu2/Rh6
o534Qso9ViYUa/x/oXnXjH4KXNg7AS6FhTKRp2sUJvcfzPx3i5tuHkms1fymiDEn0yQ6MylcPlHW
0EUim2NyCnNH9tKq63xaXZZI088o0NJG90H8+x2Y0NOZRR0HIj8eBzYpQQGkUXxwmksxZDMgTEEa
jUBAUnKBzhKbzp+DWKl/nfF0rhGYVLGKanVL6G4xjAiXyQcTEO+66nwg0WfsYm6y2cqFj4XBFQbc
ySOv8jiiMg6/JBNnrhjExHOK8PHEGQcPDAtQDG88Z+SdYRdtrRxeVtzKDNuVluK7kS8Nt7RA+UhW
AsyRpnCM3RJN0wcrARTPVTgBPyfCwL3T/4C7LGJ7gn757FLKa8/gDX2HNK9DOtrsFhLHQSb+iEVu
Y8iyUtLUSdhsTJNa7JImZ6bPL62Y2fWrj6PIBhVgE8awDj4SrGfqire4vycvmhfLYeuAwz/gxngQ
wywIZl5/6LtkYr8pfDHJ5IaPdnbMLuGE59Jj+wDAVmrYoe+j14nffLz2AU3VO02PkPwwIcxlga/0
zNNyd9LuwMRBhmM694z54zW7YbzrR+sMaOhUIvQEUI/Pki6tckuFpNJZDDHjYuhb9JIXpjQPAhuV
sN7uHcEZVbxL6pFr05LEQbCfgjdDALIYvBzEfDGhKaR1xdDCg40+lKOXjErSoaOi/0/Kj+jVOQTY
rHD9XDwMwwSqZPzUXQhg+cFotUS9G0O82WRWeCuIxe2rwpQl8zkbOkeoXu+TxBeuBQygeyKTFSI/
o2xLrM34pyACG11U7KYTr4CxEaXaHWDwgTM5ViJ2Cvu6/5ohi+jipHoNtPIP1ML1oDUMYR2uFQaa
DJa71mPX7O9Nf7s3jG4/cox/55lMuX9fq6R+UjSYXclseem4AOgAqgqdp/GzYpkac5bdIgF6LaX2
ytuCkUuuAWKVZ7RgZcVjvZPrWqNWXw3VGjFkNwA0T5T6C4P42Jy8f6QXL2iBs/ossDHnzvvRSInh
6nOemrw3bbxLHjWydrOhbvJjLoFTf+eb4Hv2AsOItlA5kpcIAM5w65h06EUTunXLWzrCble5ILQR
9Cy1sLbWcfDtCkkCiIu/UnU4Jk9f4/B6KaWoiJj48TjySYtiO6FlrKK2owhLi1iozRRfclQBio5N
6JwMn6fzm4/gYsncOiGQ55vdMeZHIimdcVkSLXtobNMHVq8okGYCdcHDNyeTl5PpS9f0Sgz7F2d0
b+lTIgqkZznFn0qpYXMbhO76GBfT9gmN47GlRYzXaSC2MZI337D2oiF5+xaFigUBnCgi7VEtSLyi
NEjQMs2Q2KLpPWfiJT7SGCgz04n38G+utCPKxqzKj4PJEFL66o8rr8iGh9/xaQ9PTIXFOtvKBNPA
asEnKsiu3lv4cJd1HyKcAXjCyHKrbBUypq0Xrcw5gVX67SVMTZ9QtNuZgKmr1oKL3N7Sx8bGKV7O
Znc6qnTyDrAKdxQbYkqjdyve7WaZZcfVk5Fvm3WExqs+qW81OqAPmZHi7SGtyE7B1n8aRGw7BIaz
Itm4e7EdxwGX2fEFLp1Mp+65X9ZTToVDFILJxIqbuQTpp4ILPyBf/IS+gWa3ZvlMTNu9AazFtkNv
PeIaC/SL+ypdbJCo1Mvn3vW1NI+z814y+3qeq/10igp1sHLLui0UXQTbukh1I/r3Qs+SGalO8dEs
Z3mnwrYYkeKeVFdTJkdxdaJ8bpiG5imAoryXBHkVxBfB+fpK2P35FyNlhGVoQGv08eyisnOKk2u+
UIWme9KOcOdiR8h/Mct0B9n3Ix41okRfW/W0O9MnCEtqFz+KuDHq3x79xwJk0ppQ44WsnP7FkdYi
NUXi+QxrpnsNyV+RlVYpBYEL/1HeAJvYhbXGU5ZocW6sYYCPM5NljkhZdUFNtHFjykocFkmMIkAU
ipO6n8veDu2NzLiDBQnLbwpH41VVFUTF8kUIhWTStP/HNvCePuZ8C5rujo4wkJEeN24YzvStNJnM
65hEH7ims6SFRNXrLOWZTbZ+lqWVBZ/q6SYj68AbXiXDWZ75jpwcQNtfeAaq0fchU459zVnJAn0m
+hAS1zhTZiDxU9LBhX9BpXbgr5kWKvYWCZ9vkhiMwNRbqcuwaWl/V3gnxnjjK4JUV3SWcOEScd+I
gdADFfRRm28tl7neZGjbZO2RDV3k8w+pvy1QNGYYRBH4c1OLFy0TILB61am4QwgHRIiJTGYen7Wx
F1YJEAiGhr7mc9kyoewdWIjU2OvGtOspWL+oVoHpaUfxct+YZ4rgy4Ne2sl5N+ElRx5m52I23R9W
4AkG6Ylrovv4q4TSfC/Bv/bgljn+aklhpOZKuZhOBf3k4APFu2reU7b/OXPheAwyXbBrlJUExaET
1P1TR5allmvc/dyXcUCWPlz9fzY3Stp8VPZPL8yEyF1cS6JhEIfINT6dy/uPBPcg7Czl16pg0LGV
2ApunxZb/8kEYsSGuy9Lzvk8C/3wg7fahCjDsQl+jcPUvcm4Cx8o7Lj1zczYVQkTpYCJJo/oO6il
JxqKFJaZZYa4YbxwF+adqh8KPrAIHvB9JPayqutQc2kko+T5SKUAhksFgYvOl/G3A0Rn/Tq/8qFZ
zXuqOyP0vYeu8BSvvBsmvH8Ma+8Ili5Ie/SPo+9HvK/crRx3UaBQ9++xooRRAUx1cOeh78BxmhT/
Ln9i/BNzAoD3j2o0S4rWuo3KedacsFFoqlPrEf/snAfMi8LlBA18zKKR8GiqfSOIBlROA1soZsoD
7kpEUwzPtvvxoX/HlpFjYIhPtCtUpc0GaayEq90zedwfG1U9tSuMWCPk0MDm524Ab5sdzQvjCMav
jUQYTa+x5/p6m9WWB3l+0D289iEJGC2hb5iAdaYFp5oGR8Zb4ZStnzmTiiCOKs6SPKCXq/bLfVsw
HH9BIi2J6xwkPgEqgcblNBaO7gEYkwXJTnRcdl2G3FMVSeLJ9Bw1WPTH2p2mRRMnoFkhu/BZDzHF
d+tf2f87e7QMqQeDAM/T7SS5tZ3L0ORIG11Yoc4tIQOjpTlV+nk6XH3avT6NIvIFy8DJfIcsCnUs
GEr55uAb0kdyXglCV9Aq3sepCVBH3BcFD4xZ3cps9qStdfuTUAL0F2STProAziymM0dpV6/ss4md
OBISqQD5Kn17c4ss7AyeezPVPWf7D4yZJRUtoRWzR6wBt2rDbwYGDLfBkqRhUQfTsW+rI8YxIDhs
3vfM6TvvrOC9il8EmbzxoN6SOQDMDEG3MrDAK4zhus3oRbJE7XCKASU4TKGHmfEPrLuLLvISWF1O
O5Mbp/zK1OqUFi16KGJ3xWaAsJl7XvuweYUViNCB3gheUo+KPIK46+7fvSThwn+T2l9yA+xqh7sn
rT8AozNsAjckk7RKRiIXV0tWM1pMZgQhcUSnRuNecOR1C1cVtKkLDFQ4XeYxrQD/Y1heeOPgbxqr
kdrVrhUYrN+cHvPyParppDB3aXoJ2+STFzdHDqKDRNfgOeGiItHLppyicpG/3b7kVsHlzfJ94FMy
QIm7NGso+EIOdBQqj061Vuevu5ApEeKdPk1AdMG2GjjlMYusPEUweVgtoVjKO4MDlRQ1jmw0973g
no/KOj1yDz2+Y31NG3dS7+bjLksKwGiEu8sxisB0ch+VfJfQzVAZ26nOtDcQ8HHOsR83IHd9ZDdv
xNHEOnhyciL6vqRWJOAuRdtWUXViNO0b0dhse5Mephl81NmLgSzC7GdXspNjiHC80Vt+4wR4moEa
gZZZCEn6A43Gjb3uRY3JuWDm0lBssc/aTAQIgOcBk5RZ7VFuPVEZxt+k5hemlfYMEWjtqrOscyGh
YFupuz3CfJUIEzej4+YDvzoeWSjwT3p/VJOcNkScBPOUmRCaSyLOLG43oq0raEygiRWZFNhK47BE
+jbAz7yetGbVRgLo9ZGwwG7779Kr6wwr//IYWgw/6G2WM6vH46iHHqu8SgkoDaZFEuBsi3s5NsAa
7+r9tunPjP8k7Anw7A8f3DP6I9g4yUf8HchVKT7akkvNCUHSYpUMPp7vKMOKVz88TiitN0qcvThd
IXoFaZeAcdrpZtHVGWQBK6ojrl2uAUrjgauLQ0egcCz2/AEAIMCRe0RGeQfxfFgsHvBAtCA+FsLE
4YhQ5ScdBShfXtyf16duBzgbzr85iuu+vvhZ/wZrbfSoZh2wvh0TwO1B3VYhsF76OIBHjge7fTJw
XBPSLz0G/kiZ1y1fAE5nk7e8yA9UwLcOQISUom5O3cDdPlvnRKiEF6hOoMBl7FTdSyYlVnfgEXEP
sbowCSgC/gOz5qHl/XoleJNy0cl4X8rDJSZC+kTQL2a6ZjDBxi1H2SGZ7qrrdk6jkN4d3kMvDVtO
5gEGqeiAbhWxtz54gZJB/p/ZymgPoxRaRJp5vOTNNqbSI+dTStWZhwtWWh6DTBtvD87Wx4EgaLBd
vOIpC0n6j6XhapsvrnizDG2qBPWHEYTBrw+JLpnIwWEazfJoiQ6b2hMXgT8LEbcW0/eIMUpbjj2r
iCEj6xrKdvHxjdeM0yhUWEHHihKDozG1ZgbYM1vCyGfB2K9M/0dojnwhoYFGViVuPsxtkQEyxQqV
30/hgF6CLFhARLKJRDNJlc3fWHjkc+J93nedc4V+ZWXv1TcuPjfJ3P1hoDKGJzF27qdwpU2glINC
xaIvROX3tjVpP+4EW4bxGTBDy0bfbrKO9X14cGlWX71i12ugInXYIPTzTTRl7lX8y4bDaeI5e1/B
naFaEX3vEItvc+CqeIn4Zr4ysf8d/KvcERs074TQnlTUryGmFl/u9zU9vMHlSsOiz+OkZyGrODIl
MBRpZUC/oDmHIqJjQgv5UxK+67kGO+/Lxi2yQgpYTmukgfCEcHCsY+TsLPRF2LrP67FSIL+6W1oe
m2TAxGOlFfkJc1YsVWRSG5EOAbluc9bR+CHQBv5Hfx6VVKqZ3riyFiYMmmQGzOnc7JK5tXLJb30u
iAzS2pZBzOfapLCrxh1OTbOHiNnb6He6c761glhXZ5VBzFGlxde1vPEZVfbNlvjd4z6QJYcOEY+V
4kWu4Gu4yWhZjMFEqHqDm7Fxlt6PBfkvvlQP77KkLU5tit6l7Uw+Z52usBdTTQMeIyIbTCYDRtbP
eJr8aRzmOGaSG0d+TCOs+rQhMBu04m2lIkce8x9a+qwcvGrroFmHV3SZswwZte2XLXJOZDzJqwjT
cAFzEUeb9Qucrizxa4ggmXqMR4JHEVv8eM6AEqkW2T5OSKYvqM4XwoA+rMBtMJyWHh+uMpFVIt8a
aAVt8mxutQGxuk5MxoSGfPfFuA+sS2GWegBYLRS3LEQ0xBoZNTuFdRGPKhhtX45h4LrPha61Lu82
d5CWnXIb8E/SGeMbhTSUgyH7qx2tzm31L0AcZdHdX9xzZ93uFcSs9Y8rtXJ7f9pUKVgfsrUvrwwW
o17jwQD5lGI3waHGK7nILSepSOl2ytkkyE84RG+p/vGKK6O89E246UEDw9tKe9jh8/gPGwD8YZB7
j+XLLZQKAGm/jrOlcjifotAl+4s1YKu5K1AC+Bw+0iGg2mpdpFmKx4TGzqaOWmhOC7gPRKuTuO0C
Xjgk3fBuWwCHVXoLDBHiN57b2BzaydctWV/E10sEvOAuhyVNB6HeWMkum0bUp8ZxUpuP5656eXWp
gG6gOo/H5HHmWeWcpyJ5qLBdbAKs7XnOlc2+yew5kwA0/1GyLaXHjHb3HsYTc5CgfTwoKQlV1Po2
p/h1y86h1xflQIgzMp2hkd8IlKKnNe7gffNkVeuj9YcpakfmNXCf+HRu8FmLYfI/b+xka1AfTwCs
fDr7PVysVKJ1gScVZRM+NQkVrhKCRHYdx3OcVHj8/0iJDBlsk/r3kuReC9MqhwI7OYcEysFmr2sv
IxFABfJPLqKjf1F2Ecl9NyJ44YVgF5I8N+ris7FQsyhlWIcQjWPsVLLYezan/CPMjGSILmFI+D33
v0c+0gp2aAvMIx2GiLhIV8ZRY6tPdWNnoX/vF/w/5vXwb/Ts9MCZCgo5Oftf2m+zQuku4y9tsWO3
uoiF6W0ziInaq+cMziMmVgim/v1noSPdOOlIg2P56fuCdHEj87wlzVuzoAmLz5zJGNTUksL6ZiHa
tpK9Ur+R6xp4EpgZzytuqQjGOE+uGyU1Bbg6rlPW6lJfJWy2NHC0s/9i3Gg7w5ndDgnP00/DnJeA
545Qpa/dD3Znm2g9/GGlZYAI2gfCjXwmWb28kCnXFZ4cJASyjx7vrv8XQc9pLFgObZ1CGE7YVKGH
DgmpyKl4I1xm0CPNyrHUsenBrixfDyjrNWXfau6r30YGrT4UsEy+8569ZeDmCPWNfkerEK0XcOrZ
qXBUoDA+9xh0f5z0e2zoDJajoTUyGAjyUGe69MmZNExeeyk1trD4aVdiAHAFWDkem0YyfC6X8Uvp
NA9FwSCNvkxhCqECB8PTw/7L0QAQORkbKI/yGoIXgtgIVG4TGRQ4VTpP74E1O/xohvdTet2qgjJ/
oI93UD9ajZsunLH02giAzJkCj6MgF1s3iAI9UOXI6HNI2ioJIWP5wfabIMMQr+s5uf3vSSbGAM8U
+5cjcrOGqDdIsDqAtt0w+E952tvqkZkOaNNb0KkNvpOt7b9QFvCiJD78RfEOdwZ4QVkiHXuSpGBF
AeD0oYt0/SmF+Cisuggou97baEHwBHMzHrp9aiNSyb642CN+Dt+K2YSL9GLdOk0TzYsdLmj548/G
gPU/WjkNTbrE8nil4OFYm/8J92ylkfItaLUsddKZZMwEYdkH91024M+g6dn8KWJ5P3LLfClw/4fJ
5/rdqeywTHfqhU+qr8iRA52qSC7QGLD/acsF6UYMN9HsjOO0ON3/p2nT9hZcpO0v2aXDnq3btBdC
UB4GBpeaRLvgZqGwPNnRVCukU3IHjyNQPSSMFDuRivlk2llrVPxUQ4ZhjB9aTOUZUv4dgG7gFQnH
Ez0IdpOLv49JHhMI+Cv2k6CF8MgOOhrxkCMzIEd5dQs32QAImqw6PlauS/mkerkRXDRzaFdbTDhP
TlpaLrZ/RpIckZEglOxf8DMxyvZFHn+CSTWzzK7gFJ4FSDWmyyh6CpjC4+VHIWIU4O7fOnJ7kVhZ
KqBhWofENtsZWAqrUBx2eKj/RepMtq/on/4Vj3f4WOAyW6P+4/CrKNz3FfQQmt+4mYRpXPSF5Jfa
HosCV/HJKh3FfteraCRHzJyznwkR7Xbx7ZSkMIDqu8kMa4b/AoCBIe4wpz6TFcVlTNnpjbrNXj8H
P+XR2Y5gUS7XdwYOMTW76BDAoEW8Iq22e8sgQRcsyRllE3fpnDdDKLR9ffAulU7BVuykZ/yploaF
dhgYosM56YTw7qFY/7Bn9+TbkowKlQrZ9PYlL3auylvlYlJhA/PXzl4DSMJbRTy4ybq2uc6XmCbB
xTv5mm6gO+DOIrnBliO0Y8T+IFtX+gr/yO61DA2Fzb4vqSDC3lAxhrStYGXXtJy/S7KWVr9zpcPn
kJfIyOH3IVdNP5Q8ffnTzfYfNaoKvgrz5+ma0WChEtAqXhvzs4Zs9Aswg2EPCMoOAkrqBJZC637v
deXC/JxqaPtkdlaskBCeOPiHMy1+kRUTkh5mb5rfbBuCE4ZBFc5N0v6PcsmgPmr3U5LQ8tfM+H5G
eoQ9Jt5Ag27EJo7P+klMQ1MRzeSOgL+K7AwV32CxV0yUoA4O/UeTZs14L2/6WYCcFJTXYw/b/yWN
6KJ5DGgXmtmSIO4w+0oXfdrF5fzqYVmCQy5sUloe6pzJ1SfhKqTXawvQYsMjYjrUGQYLxNChSmED
lG3/c3oUxwcmRSpY7YHBLI9RbLWHM/siLcKZK+8U7JcZNNFYcuxs+54mHEtg+XgelvkrCtw7//qH
Fg8IWZQb8y1qN7l8c6YLvsJFOU8QW3mVXrt1U4cNR392NfDKGmh0XvLpaNiWXn105vcylOFYJKVF
gdE7j9kp+09pienRKyc7t//QD3LvUkiVaZcKRywnSnJ3803Q81PcUWl+T3Ad9qUjLCtMTnW4a6hw
02VhXeHvICcsZ9xNwHQxBgAV4vMf6mBVBXrRSMk/2+Bxu1qb2XUfE5lf8YQ/03iPcwC4UdSIFqZe
rp0cmvTAjJZUSEIrzPCH/3iKyqRBlfCWBwCKqMqXMLmIwWbUwqIc2V+K27AB7FDfDlCW0uuaAeLQ
kbdxdmkUiabuWUQhYUk0CZf5X11y5D1KYgGK9xPPbkvOBc0omaoD8vqf9b9CrLowx/Y37yg1s/p0
vIMYUMiZr4hIxYiWMItlx1XijrRw1ttetcXmhcbj9FFdH8+p0JJ7KioV3+zU+V549U3aYPQP2WHA
KIS9J9RyfcG0URcMkIfEzcGSvqF+fX2ZZrkSqPp9VIDljBiV35xY3DVebVPEXKtxIrCEkFwGUZZX
tEhene1MmuAmGI7j282s7qUc/JnY0cx5tKZ+h43n+85dWfk8dPrtena8aPseNZCYnfcQoPLxig6n
5b0qM3IC/bh6kbm61tmWJGjaRIAjIr8yiL37F4GStFEj8ZlbVwMCSagD7kGw5yg8Qaayt3ODBiEj
wsyo7zomfZSyUhSYiF3ZBjxICzACUMuK/1pIWwcuCbnd1CZxS1HuPj+OR+fHa+BurmvU3zKniVCw
GencAyzJ+5vQ89naRhRqt+VHSl5ketVmuACg/bVAgQVehQztIrdHAPsHdNX8yOLrV+Kle0ebIprF
UMSpm5eotnKVFmV21C0mrcsO1yRnTkxWrDDgXoHDKt+ZyFP4uPCD/2kelb2vKgaKTcVo4OUxoBi8
+RxdrH7KTw7Ep2KQtDpgDtmcvc7jwjqM/aIWQ5uWkoQT5JiD08Kti9DdSCZyYbTi3BhVs1NUnEm7
LCfJc2qBhnqjLVU3D2EcjOTluU/O+/TU5cRR4MHHay9+kpeie8Ma4S6p3Ae5L0iNIiCjNbBRr/+F
EG1ORfnQeBNjE86JLwC4q6hDv2VyQYTK0g4+0m28Jc0t7AdXtwUkJziw+lE2LlPR7rJa5R2jg31r
UCriAmaBRRga7ku0KXYJ2zIBbmjdcVU15vxK75FqpXBLv2H8RpMZv7zq8dbPZfmAwCOMqlvW0ydu
GveecCzXI7HZB+IXu/Vf3yEeB1lAC77lrUOCXThT8JyMZ3/lTt69091iPYqhfWGKPdtKvF2BwhAo
PTye8WYqEG3N7t/6+ycj1Yrb+KthQ1rK/UFjJwoPWKoxSpokTMsfXl48tHSscqT2sR5k8XK86/Wz
gsdossTHcVdHOWLc5HOdNLOoHg76M9myU2/nNfpmHeXL4KMa7NzckJbUMfHInsMbHI6DLO0r4C/b
3jFhrNkP6MmDokd7MdPw6hDwtta2En5QsjFXHCK4F2wvmiT3bPb/ikINGwTxTPLWtrnjZpps/Mym
xJgE0TEqFDISImz2U1O+aUz/7vJv781sA19wOOeCQNHGivSCbanva+3o8wZXvBeQjwjMe2dvis4A
hApJeJ+RBignXAiZ677mkJWewuNvvGYDjRbYsMvUTq+LLM4t82eaN6aMl7y8sUDji4Sxlc4CV1UU
zT1RQ7VBl8kHNRuLvCrqcWpYWsDbkj5ruwvENjiIxiscc9fabPS2n+uTs9dDjrgXnSN2wpaq3b5o
KT6fUHz/FrzZrKOUPZQHkvD6p5KlLzarin3h0cZdMBG7kaXfiN8hA2eo+2WI93h82DyUI6FYis5Y
5s356nuofjsaVwxTd7wtKUIAcRMa7Tty2zFW+zDHl+Sl2CPVjSL0pU9T2hr8fpWFpyaqaHsWPIHr
+v76ugMZlxphvjmmdxxeZRXUs2XxNZosT9FpVEmkkzPC5jRL9P5/pV395kQA5abCNpnDuRprGWEO
yD/1b4U462jtITBgc6xwvr6BD57aO5OMVVo9B3AtyK9Wc3v3Ety5Ux7L00oif/fymgGeYlNdx7eB
7ckunLo7iIMkSeJ4W7P2qQoc3g5iwaSoqUxTTlNzJIgwY3itaAM0TRUZzVPLQ9Y1qBAPDDR0YsDU
bT3ffdmxJ8xtTqnaCpruH5mrDU/NOHEHt/WxIiY84o3KEBxiuSkRWz9gvXmJ4hE+h6zhipAj9NEE
bSzB/kUZwQMn47Pu5eVfBcOyXQwwBqvTE0GzLAI/KtJ028t+2HAxTSjhcGZpFarBXo32tUfj2tQS
e/9ajluHFTv/EpMMxBdGu6AMrauJElNoS0YLsE/TSN//BWrDdtN+sav9Qiwx0e/55kGCwhK3r5Q+
cHTYo2sQZ2igcAHNAE5SAwJFXiBLnLMVUH1xfbqSa2hzG0D9NxSSTQm/mi0Mo6lNKnR2RbDGEBs9
kE5Koiw+s+BCklC3VIgkJ5lsQdHBPNgyVqQHW4jzthv+VzNMH6K9VIqHQLpMIuw/jCAgcAeLTP3c
TjfFUi2lc9JBotSSL6ol4gicdg0W6xewHa7lEEmTRxleadgF9Bhe4IcVPTaC2n3B1vUx3nfGk/zz
9qgyETH4r4YuiKpVztWkbpRbAvk0M4nrPvq7y6MpLy6KkFzooP5qOrFB47lDKe4LnN2SU336zGqZ
rixd3XEE/sfHmb7K1yBU6vIM712eTYGLeB60DiNccEHtfbPqyLDxZVO9coxd8JCdX9F83AgoJ/qT
XOIPhWjlzRfapPB5tUIN1IXvCMI0l0E64F+FWABfrdQXMi4/gsF1YYN46rwjKrFNHewzr/M2XZZj
Hep5KLBuAEo6PySOweyKZce22FTx2OSau+gvGuC4lv6YBixo6iZlN5W9/rfLxZuUkT2rBWK8RNXN
AXKcYepqzIXws2v1DxPHIEiFDmNJRmrSJfUifflBfyHSO4skurwh1zhM+3uEkkL7gyEb5zqPTL8n
LkGnGXg5G7UtjBk5SD4j+rzhoedpMWZuBDLmDoaqOp0hBFXf2P/WacEaoatu4TkEE9bY3FLtZCWf
YhaKAvjZM1geuIhbbT00xBz7LhewPkNE8R8cgjp5sy+Nc2l11co88xv0OQSfiexTXb1yEf8Ut4nr
GEnS3F5+OW2WxGYHAhxRdOnezJMOesBkuEH0zsdiUOzQLPHK66dPB4x/sDroFxdW++6gKvgBgGZ5
j7PvaIBbMTpwp9VF1vK7Up8anqpq5se7VwKT7rtngQM1fo0y113DgCctgY17pqtXbfve3JW4Z7l4
44uE2GzJSkUx5X+mX67R5p39X0HNpqruIPTaTdLPezIRBLh884iRFU3ZXYs8zjWVh7WsxoehrANt
J7GmsJs1/liUueTYfKpCoQVTyX7tjPBgqodR7RyT1mWMCPIxKKhzUYjJuN+KYNMpHgO9JIeTs2bJ
soz00Rejysmz6Jyzhj25+U0cLtXLW5DvGU652TqyK6Jb+1t7ax4FwVpZesNTzi/fTB32F05muedw
WPTdINqyGMPbCSV9VQwdhaW7oyTJuvcrHhUN/mbP4KJVqkXvDrPQX3Za+w/FrvGprOtC/vjek+zS
Fvqt792jC+a7g35aYnOGhkCd6B/qd7dGuqfE3i6un5pFAbIm6AHXUVg7pWtYPnBSF33zAOb5PgmP
KwPXCfCjXl8rH20022x09FG8TrsPEiJ77EicORitrOPKBMB3bybxKZbNgLnKT/jSPoyk5oSdNwHA
7AXnmGrdcjNcUOweH1y8Zk4uhtd+t6GP0urQ1BPugVnCi6+iJJ8JWU1XT8ygafsAv423HnyMuGeS
tCZBDqBuLaEfujU6/kZwZiP5eRm+rjBfmDrh3jArrHvEv9AwsGbaqv7gX46hXJQNIhJHbHlKD9+f
0FO4Uo7ZMJYrsN/MOgjQET5paqVze01tALjJdnhv2mkXpl4JqiFdJ18UD4iSkJpMbzN+0LaNqQEg
JlvqsVK5HwV5fxiWnLw2gA4jA3yt8KwrXp9PeeKS+QByqUvgk/2HeVxK9zlsRtBqOrPZsR7XlzGw
LGQDSlQhM6L56KPeBnop6Qerlzc9IXNE1DFW6RQoamd8RW6S7LpRWQqY2oPO++Np35akztL8nYR8
FBMZrYOlqXT/pXFLzTIF9OLmmxBwNoQYoQbGUi0ehw2VtxEF7VHliATbo3go+jITQ0IkyRyZbSwm
1yZsDha8gLzxCFncwouhQsQ0aL6ia1GFTBgYyJNBnM2uqk+WC6vl9W99tlOG5hZmcIcsNHPlwgHH
AAPY6HTLHF2WWBUd9geqzbD+/Zumnzj7r9cgRoUPup9V6bjvtX/t1aPA22fGX7nuqBqQPBZ6sA2r
Ae3T7fJ/NucicG1Fyjl/pxCN3YLjUrClz3P0gkB58OLSrriI7df3JwiMxQFjdmHcxzF5FdtIbLhf
3EcOpQuRK8EfNsjaXGya1exBrtsXsCTS9T0P10th888S5P1l5zYRg29BnXLcJPawtZN7qdgeU04X
1WK0BVEEhtYSvgkijGfOxvbV9rXA0PToTqcyLMpi/ddWqBS+33UzoT4uOq6UjZxvthDJHt5INIjX
hO7NMt85HS+Uc4neWOqknwDk1hWulfyZlelNOSpBBx2pD1dUdiqlIC1nFVZo7s3F3gFvixJa+Wyd
fvWLFE+DboZv1ssN7yEaoPHv6fFV4StLzxjBV/hx79uNzwAQ+9D7COtdug9F7HgvDe23Yc6ihjIF
RGa5kEI9zOwf26xS/lBpUtoiTrOjANU6NhVu5zxQD2awEAOMed0k76jZMVGntYdbrI8pSZnB6nec
kDbOXLy5Nsx9mTtbKXJ+G4KvTiMNGtEEP8jObofaHGHBUBrZ7z50O00AQF+KLwfWpoP/nfDNXl02
CYqs7YaP/8SNVRyxVRvLaUUJmtCIXSAM/By/s93BTplBet88ImFtC4ktoEnhHrxRoD88xwANBgHh
04OxymVaOOSuvNfsFrU6MrO8uVGbNQ+fRfxVXunBG1ll2lAXiPoB33wKy/3Mxd/Jy1cwYT4FrCCv
uSvjUhTlyF07p3NtjNuC/lXfNK+XmiUjyA+fQ5S6PSSUl4AtAuJEjW5sT27MKZGbbno00N9cRtsQ
FUK10PPPzP4EvzpIokwMJrFx67NR44fRDAjuFtKr3A6cMj5hgb2ypPre5MNANRA9w/lFlQOTOJhy
4EAsHp2rX030U0YqHjrlpjj3UYfper2QGApltDpAhzxcLQm+AwyFjx3686VphkPzun8OZ66nGnCe
J5Jx6TmbEt8kvL5HzIGyChjjDw2SymcRyrJzyD2FeoE8kYEzmzEvxAybdIi6wtinu61vje3FWej/
CCFFGcrPMSx/jHJoN6Xx451DPVlOElOKzN/OGpJM1MNrvg0c6Jh2J+rBynSCxECRohelS6Q0p3Ce
Bylfrmi0RXPvyvyW2vZhihbu1hDWhqIQCIP4mkJ0x86bjYRpTHf8sA2siSlpA+LPiZwaNP2BHAUS
nkx0EZQ8MVI8X2Jpa8bXXlcUjQrcbKIfU3EkRJAPR7s81xGHxDd0h9bJW2PWtpl9VDv2ZoTcgc6H
uiQN800a45uETNwZUu0Qp7Ld0tqw3ZHq97EfsGvhtUGFmcvFas7Kgl3og5bqH52m2R5d/79uBpbF
D3fK4DQv+Vm/yOLOQ5Gcg3dgHBf25jr84YLIkM0jv8EZsbkicz7MEJjI56i/j2gL8k7B/AhFhxWW
e0iRvdj5E0OKEMY5aMps8Oq1KFOiSQ/lkdZCCJdTCoqTp2rCp/6HOHdiLX2Usx2TojNpFty0jJhM
mrm5i51EDUeVb5V8qFmlCnAJO9gCLFxxTC+QsWrAUngZ3JLkDzF4PiUW/AniDCVYu+QnwpSKYPJL
Gq6z5E6UEiKEZXddpH+1B6alpWrNwWgb3MuuGTBZVe4xP5/d9nlh1r5laFqLRVIGTtB/hVa+lZd8
b1WtbDitbivgomkSbFe1fpRfpTpQ31jebDpfoh+qrA3KBPY0RsLq1jqHUeQH0SmRs+dYhHbQitac
LO29yCpVv5fK/6FBUnfThiwXK/4taBljJwCtVLXhDloamy1gT+qqEc7PkcDkRcjnPWC55YPTWda9
CTUy/2U/zAcmAAzQJP7B1mkBPmF5Dbs18/B+4JAxDYVnbNEnyQYfsra5yhxso9qzucLP2d2sJ7Xx
nG3vmguJkNQ2tpLNG6wPc2xfBhdJutuQ/cOEjrIGEeYANmax//UPglS5PHVGr3AppmBlIoZixauw
2XVpp0EQq5XilK6iy1F36nwNFg/hhwjqk5Ldpe6s75LGDiA0xWg6BeEmJEcmd8Yuopl+ZdzUug5e
dUUTv8kXAPwgLnRifdxVrHN/AbWhW6XdbIrfteWiphJ0900NGR72OWx7AmkZScbjWARZ0+/iaYbF
Qi5PlT+jLx81Ky0aAlTsczuw4AkSirTYj+5dybR7wMu66UFf0e+ckxi6IGOo6wl9IYES0ix44hbE
kwkZkaIeERcEmNcem9ZdIj5BkjM89ofyGWXssb6s+vvFY1LJa3JD3xSqnIncBIz1JuDZwTgPVkGA
xUsujvNnIOFWvbYjhsuGA2xFnrnIi1i4L+CXEK/nVZYIrtiy79B33lf4J1Sss4/wiaSOE/Vi54ks
OJz8mAE5AJGZkKhJDPlu36HTTNtDIy6n9kHw1O1SkPDItt6Cuw19v+sXaTwXVE9mBmU/v58fhnCG
zXQhoziCycJ/XiLbqxsM3cE5QQK7pA6shjdlvin2zDYgT/umJ8HZPmDXS/Iy6xphImtOTDkDknco
YBxzO7qPDMqSkqFjtxl+w/vQwH2AFXej6Xp5CclNdX3ybRVnSynVHJ2DykcBA/1xc0eH7XFzVtVY
H/FePACJV87YP4t9FrQcq0LUs1hJk8IoHi+FdSqrz0w9yyCDI4O9YWp/yv/EcZZS1lF3BG7SRB8K
li4KXBIENteArrTK4pjicbISZgd+XWN2VAOaX5njpG//YsL0to9kOhAKVnokYRJ1wVKyu8nUUsOt
0q9le2DN1+YaTj334+4bBeMZkWYEEvLzxPZ+F0CmnYKgyng84x2iWJvfhyJzkWOFONUf+cO5WjPJ
7Q+1xN375+zk4HG9YmpRsTG7j5bBkCqDKEeswRFvwzzPx8hSmZTuLdPZZ8lpXzmbPoZlaaS+G939
MSgVT4y4UJVnYNLfmlu54P/dxyOYgmk1hAIlJhxbSoUALz8O0w9OOkzIkvzNwjA9bUA6KKMQhaC7
tRPnDgzvyDO/zq0eG/mdp/WKorJBlwbOw/UjU1rUlCLyDi8AOxrEsbVGcE+KEYBy4CIJf8XnXfRb
cjnADV0yHQZAsdMpTOqhuRMaHF8yBdu+6vbdWJIqWC3dx54kdWQRw/0vxAhG+wMYXXoOv+SnU/jd
nIe4F9c0UiwuSNXvAHGO2bLphbroSMjZI61xvfANnD+WaUc4NwGb36ixWxKXh0zRA8ZJhk0/UEzW
07EGYHsi9r/JIHWPfTXSYNzVmvKFBFbWMr/yzDa+tztE4/i9rSOpNdkZYXhp9jilgBLhPyhAqgKL
EIikit63i8PbE04iVac3f0yw8sGOpHr34JOdh0VWSICR8fCaHyaCBoRMiNx0J17nf1FGi1miNVZ0
knF0M0hiJt7onBOU5vwYYsBhfSRSHHGQRq4uy4HSXFLZywn6WyJ1kX+4QbcAI3A9G/xuUnQKFsze
R+huQbbzpfQPoj05oDSiN03aYGCNS2Po9R/VQzwPuxRkqNz889oQ/aXaseHig0+85iLXVe6FS3BX
NGMubgkmq+VZE/jB+ISSWjT7DEQ591V7FReh76hFlJdchr2pjWUGCC1V6+OcGLm+jedRjYh6jbQQ
xnWFiB2BzRU/NmF515tYabL2YzLh1VaY6ur+JHOsuKN1DNbKC9EYGI5QfWhoBghYSvZqqcloMSK1
KQEoRE5erbOEg7sDjiGugQPRPwBeLAnSfBBHXfE/qjs1d2QWT+SIm5pg6WzbMVnBQ3OtTtpx87+S
ivS0u5VhGW8zYOcDrPSab9aVzNr1oTiEEcoXZsGigyDNhbFSP0CJ9Qwe9ad7d11SJ0OR7LbiyL1A
ZrzAlSqdk/AOiPoFLGmebvEapz5WUQsSv0y9dW2gFnhHFrSW9JPQT4NHgbvlFSXnfv9qIP06Kb+X
X+tbJi1q8fVM++vvgdFMT4g3UthSBDuKoVgQd4nyvssRs7Gltwmt4XKL0glimdlmBuba6XCggB02
H8sjqlHckD/YK/iQorLanKESaG4ZTiK2pPWNayunsUrSEJofU1tV2HDZigasRkMMP5012m9wC6gE
XBCWu5UMwrUHT97PeYmxsy8sT+N7FkrbUaBB0YzENt9JYGQ+211A6FDJ/eplWsrhgmSswFcXVJ06
+tG2eKS0TSk3It/granwAbgt3fmoB9zQfUipCe0IOJisEItKctUUdENoPwclnthtb73CjmWnhQ/7
NqcZGLBLjxbKod86sCo0P4LFS2j0VFgpI8cAktfbpbePJB21YKtSDNkB2xFeh+Ng9h9UuEbKx2m3
uo9wf5g3KzlWAhrKOptzNYYJ1sXbaznkRudW1r6GN5DAYH0bpngpt9jvcXUtGLOtJU1H15yMw63s
cxDAlS4tz2g4Dzt1ES35SdCkhgJL22TQMqO7RNrhfrxhTH+7Uv/3gnBpQuZSKP/KxRU+wIKHmvVz
ifW5eoRzG92UUnumInNz93GIQYRIwNtOI6v83196AOppra7m8IZMk0r7jTkl++AJ3mJpDbrYrPVR
kfYFtfna0Gs3WGyJ3OhNP9wMZZjbzIbyMqf1xnSAVDSPGHttTIACexdtMG6zSUH9JioJAKCLE7Wj
LazUYuWLSKxky7Gv9RDRc1mcWTJo6kMZ/vbb/eFHxfs8nPRsN5vlDjioH78xp1SJAA2PtfmCgomy
sliouolLl8HxYzvHEneHORYp8Cc2dBTLAbup6gSii2660ImCGVno7gN6iGVn6MXa27fjLhSw88Ro
0zPMGwWrcJItoPy84+AZnhciL6hw2IwHAOuHcYtB0RSNpGrwmUHA9/tK1u8w3hJ/bV7LQgrp8SQY
zSYIDjOQy8H04szNNV9hSz6297ojQPimkW2nlSYEfjSH6/z51gB6KkudOr8QP6kZnZctbg/Tz18h
c3IHuhr/vobODoUHZ8zSTwIS2phxhxQS1fSZ0bHWIVV/fV6JRVfQi5O/uCGz9wwb/gJUDC90OK68
4s38n8/AzQwu0zKPzegM9qJFQCOLnsPfLbJ7LqTt2oNV9hq2Mztkyw17OirvL8jlPBszOc3ysy3A
owOZgB/me/cwFs4twM9Q/hIZSRQ0tpJq0z2qawIl/jfwCx2d0IGpV4fwaLeaUociRRbVBuObCQVY
cjsK0GSmo0TmPwuzhHa5/yxzuoF2839qtZ9lAJpVh5Xl8+dBOj87XCKg9WoKOl94P0gyFUHhBMeS
Okk+2zctOeHDBF4BcnVQuVk0hIF873aGT43duTAzD9PH5l+Py8w/nzciQrwLcB98JdPjSga0/2BT
59jP+rCtYb9GMeXt6Ky+t0Z4J9nEsAzVKAlyjpLGBbLqCZ3w4FHRk0vZMJqiPpQMC98xR4gFtTm/
TfUAp8SsiD9XsysQqXkHITdgG7pUNcmnvr48fP19LnE18ZJxx9kSf+vWAyCc7m/VEHTrePuBUuNe
F8B2z3yctrbnJiNu8oUD9Pybah7Vi40bZeKoV1H91ZrrQ0HGL3PkKKhc+DSmCq2opp0d+1TUk73W
Tzleac+gFnbXqo//J1WNj2+BDv/NTtzHpYvOTslxfL0t5OokXrqd66XyEaLTBFvpE4IZbjiMSf0P
jUS42mFI2ND/FH0mT8Gpy4+k+BSUxQUb2S5ZclXkJVsFZjzR204iKkXOR6d0HCz9XErdPu4sGEO7
n7g067x86cr6SsOB+T1FyTJKFBK5A0iVWuSMGIkD210jyxpCgwvH0bKXDFaiRBunyq3PquteMN16
UNkNBVb2IjA+k7FdpFyBM+UmoaQn06N3W3G1qfCjBc8iRA0zMr1qGyPxXA42zuLlg6Rg/OxF3ewV
UttdNoLkXmTk5VSp1llu22K0EpEk0xKVc9/8/pVi5USyD40XxRgu4QBkhSdjbmV5A6hkMpwfJUct
UjTnKAxJV6XkeamLy/3zXcGE7qoZUn0tq4xqIaX7bxYBwI2gbB2HehRKKwGPVSPbVIVNYkBPj/n3
cGl/xGE0KXgTTeUyUKsPdeqDeg5+cuX+n4ULFSNkvCnO8k6K0Moh7YZ/K43wulPTwOpyjjznd3cA
4C4EvnQnd5J33cWqCsYUT/KCezdWEFRTPkRaIHpC+RpeXD7CsUWqKY2atVLXm7wlOX1SaTRL3Pfm
3IkdYtamyJ4phgS90WqEuWeUBYLoJgs+wTSB7pgohz9TC6aYiuePfm/rtpStTmKaX1rsHT0lBAiJ
Cy0Z7MrYmU7DYMoBxDDK3UZdBBwUwXyEjuoMsCo0gvd6OeMk54lJgBFLJ5XGCMSz7RydcR5A0t17
SDJnxVUgOKLsF+5Z5rp9UbiMUY+OxGUgQ0j2SpizYeArHSiBx3DxJuMyRJhn7eaKDB3OpSuBJ/Ey
l/Or0D88Do6Eoo1GKe6kvOqOUYpTfiDDo712KQMaBSe/B1So297++aE0Sh+638BTCpYVmPW8PX/i
3IqTm5A8tvu9YhfMTSBFpZYRTh+1huvRoHatoyQN6IEDnu372HllLFw+yccy7a7YsBBVjC/NSX5y
zGkoaJhmRVBtbCtYP7NF8TyOl21pfTSZGz2SzDfCyySbnvZgw3czCNuaToNN+qjML/B/pRX144Ls
DRvgbzOg+M/dd4iWFn9zOo65SKkZ6U1IQBztFOJXME5VNY9qJrAm959hC+VuB1qKe5UytIZzsVHG
sY0UvnQ5M0jIhyB/sb845UKcZOn6flXECeG+xt9iWwTrlbkGPGZAtsALAs5MoL3p9CSIyYyTjxXR
fdWTuGfkMNkiGNU4zrgYM2VbX0ju1tgGSBE97yuVedARLHmA5aeZ+Jgj4qHziNTh/oWIv88NzYNd
jHG2PKpV+6AMmzBkzPEQAyk0tFMLTxTttgGHiEX3fGBBJY/dC9K9+z0qPrVhkEnNIcO1LUIhioMI
LABXrJDa5RyQZQGX9eiov5RUAZUeL9InR76WLSz1SMnc6jKRq4g98fqbFiB6RAztX0s2Dwo65+Gf
o4Tewo4xolexgpgbRySZlSGw1TYml9Fhw3JId54WI/x26uP3gi8IIZG2umMDO+XF2tPA9gzbz9HR
zURGGqo8ZQrLhfyUFs9bmfTG9/BJM/LLNEXvSZSWK/EEyqkQ7J+Jka6UktF9/7XjBu7crCNkkMzH
+B0XOO+iImOrI5w9v6d9NS9PCGeOhpLX4VyHOZwIge8OTd6KiokgqDeMDoO85HJB909Ztp1tAjpn
A9UBu6BnGcXEIclauVjBOdeQt6tnZjVbHB6tNTj8A/RnwE0E9Kv/dDSr0+TOVx3RCKpDnj8Oti43
1mcmNxXOrJYjWOh4lHsV7lhmDgSzBROQIIyA1k2wqPKrUjQSi9OoSWFC6NDoaT6jMYjey+Iydr9s
lJqdEO8A3w5xGTiEbhKe2EYM7F4Br1jpGxnjayTI/SGO7HTJle8nsP2a+pkt3d36O3jDfZtA1Ol1
dmqdeR9PT+AsLxAlfmhEJuO9eE7xFbwhO5otvq9A23HLVcWUAcbJYz0KU118XK83hzT6W+dAZg+C
A0KHQG158Okr1qmCmmlmIJHdtst0Z7oe+l38+2yv/hdpY5WQZdyPDTNCOAN7/8NasBffOwbJoU+u
/Zx6cx+nCqib9v90pZEXyUQbksA3kMAxacj9pOYjZm7xXW21f3HSd+QdXivXa7TiwKmTzXSsT6Xv
y8RSbnGfZATZKN8eFPNyEOd6qJgLLE60d/FBkM0pvG2iuHnFtipA7lFFlFq6x9mFF4Cmmq1I0Zds
5ogzd9utmYWqf/ZaVU63/rb5+U6CNSCXuaSsdK5hMCzvFG1yYl3vpNE/AwGn7JakvrUhkQX9DHe4
SX1/zaRn36TmHLjLtouinV6IymCfsLxkkjP7ub4yJuzwCpkQCYZrxGLls706fqXrDkN/nfJ4X2kB
BFHc0GMaGS3J2mBduUMmOjrwuPZUkFf7EQz2/YO8UfcyVezeedkyQo/3Tuh1O/ezTWoOmCE/iwc1
fTQAFsr/J+v3IfnOriprZvo2bCADXkQgiXSKw7rEp86TlUO39UxiqYokuc0pyvZIuYXBtjSPPED0
TonpEHB5VamPYF4AhnS7LzwaG7UZ28obWtIvPw4CZRNyxaeBaMLUtt3YpA9m7AY9ZG9DHHg9TD4D
cVkc8h+MTBsGpXTe5TR4JtierxthRcOl1g9rCGYd1P9z9uh/gwnB/HgClFk1SjpH9RX5WyXFdHNa
LrHRM4/2T344xZwcC6fM73FUjOSRpIQPEGiYvFuaFKC6ypf6ri8OnVndrcMm+IFG6Wv2yErVVqV0
MBEKiffKWeff8KojmgVuSMkmLmwNwtD01ggXiKmncr39s++wN0vquAwwVzJssob1krEzRIXH3lBi
kHmShEBamxXF3rysugYKnQP/+53+COrj4fWbtDVO7uyMNYAxn0CLOU/aSGXqffaCnZ1Bi4PyB/jW
Z/ABmvwuXjUO295YJKinX9hw+2zYlLgG52FNVWtuoedT0GDdBSxNBsy6cDffgXXjXvMJOJ6SCC5C
x3u5pW28DgUTs7Xnzbq85b8+ZNlMvg/mLMsgnyIlZdVPTFPipMtosCvcOwH3oqz1fh6AILmfJvPP
TfWROir3WLbFvYpc7DIH0QZCR4pYRpKV1ZpATy5IZJBh1EFAihATWDonuNtuju2hXu0OOWDZKk7Q
5EDRK8qd15IQTas0e3j0oVNOklyZKhqxo7lReyfuS1i7LFKOupKVytljhW34atSmChfsUkkjP18o
mx/bA7GcakClHY/1n8Hp9ZFmNcDrcIqTGKIfzY88mT7QDKc+r0x3Ll0yegh1nnVZy/HA+IVekAo1
adw5S59VAL4dz0cKzvoryuYkEF+RDmZq1+dF9xVqJKvfN5sa63GxwzCEfyDU+s9j/0FiGlfakPdL
7BWOTgi70vtzKs0tVWEbCYrIkLfW/u1+8RB/nVCJNea1ul3r/+drNrHEognjDEpCBtM7xIHCgqmG
0SkHrjU9GLA9YleqpwJbSbZGx44R8K7fT+IOqRfQTCGcf87efXqMVVa8rPRc0eAF6cV5Px7sUHV9
F5gM+N0lStQ4xwhADrwtVXqGkp6RsMrkOTLLwqLJAhQcZTFLjQC6y9rWwwyZFQdxuCj7zb5D0fD5
Rz+wow67mRwxD7MEgJ8SPPtYSOsOWG7rbsjsRmB4JA/ZMcqPhOJtrUSjn2PHRtXunqGayI1jGjgh
KoCtzR8XRdGc4QMJzLFjj5YgwJYBI1sjej265pc02g+/bAsJW2E5mYamXirP8Wu3kE1tLi6oDVRP
z41HP9JWDrzRxQluJMDTxgW/lT0CQY29xpxN3gS0pKL1/Yvalj69uEaa0YUOzy3mBZ3uitS9DmwX
KU51G2TM7Flcdj2KbTuMi+eWLD3CBQI/8eu6DU1N8xFUEBkbKKAtBeTlifP/uYudTQkkM1jrVPjB
TuvE5LHppvr5cjhoY9V9+frBremjjjMTPQ2ZHH3MIwQZe4p552RtwxtvzesC5M1QaXdCwDrdQJyU
oy+rxyhrDQwod/IkOlADii9R3cn6QOUF9N03MLtARQld0QqO8yf5JFcFN0ZudbzzQzzUhvajq1h0
+QdBoSxXYfezK16AHprFtm4gMhUXY3Hoc7wNo6dFavTXnx7O8fLCERjtKUoIsX3SDq0ya9/FO7HB
XoIytL3gGZhXC321lKMlg+5mcEM6RV9R+uBwzEkY/oQBXSeHMFNGp2Ra1/JJQf23Bnx9UL9cOCYt
qggnQNgpi9t6ywYXVulZMvcqbnBfsaZ0NkVcp92VdWJcQc+0iDI1EtY5dUQSSKcw35TO8s+k1VTP
f1RTatrCv+80Mz5JHUaUqwe0UdmVjrOlnS5rhHcbe6lx9fOL6oyXQA5C5tG+aq5Cybj8rRdFa0HX
5tnuQ8CAbVznF7kKe14jq4UwFnEA41CHPO3goaxmfhL5OyPpIFdHm2QS91B71KzaKLixmoyMUZ3w
kmAup4BVzHVCmlV+wDQckJDlgVP2ZNaBkCoiX7EpLeB9H3NWSV7fwghJQPYcEnsANP4sMI49hDYP
6fLYncx6oRWKKfvIJ9HCS+S3y6nc1w44tkboOjYGTrrabl8xWa5UIV90Y2qgnEoAEtd8+D27omIi
2CbLr/y/cDTlaURoFzAmOOwe7vRltwIiX8/RuPpFGoYbiXCwp04qeqWL0fomSurBppQEwzzVWdQG
tQrFGUexRqbBffMM/EiNQrI47kMh252e3p01GHUCvkQPc2Nx1qVly1NqYqFV0Bl65D6rs0fXYvWe
ML+55AqoTtADucuqHz+sdZQIksY1nNOxE/cTP+sqmpPq1Mq6EZkYK0dceApbFR53Jvp8tgT1XeAf
gZh342vyxolIb8MrTHgdD5XcVvWL6aylElFDaSsVm941K5e7RINj34+bFXklpSVl1SMqn/016vta
RG0L09XhNVOgJAsbntQtd7AW0JfXzewLpNub17jTX0UMgg3D5CWRWWDkpqEJTd4QoBgIXIqoCr13
srERmZYvAYJzOpPF+w1yJd5qSm0tzFJvkz909Z8L/ViEPC8sBUkw4ABbdxay2PCmIJaeHSmG7gbf
Ek1w8W9DhoytPwodEEZC6p6LvZrTQFxUViQuZ0Te9vugytydyT3+VV9uEOOyLe/t4yPWe7BaSalK
D7U3bRdrXUHR4KIr3gAs9EYk75iYcvre2Wh7MjUxq9qpMuEpvzyv5J0AeisMToZLAZwVw15fXEkR
CMMIQmLiDznnIlIqV45/usem4ofdzpGt3WKBxjSC27xA5ge1wo5u+adZIC6cR72EDicz5IEmGJoD
J9zCw4DNQJu/XvOpK7GhxV+1Uxp4IE61yEquPf519x0CmglTF0U2kuMdpmkeJGtjFcvyjWpCLGI5
6NRfUkXLMdxLq52YGFCIGfAznQvMsw6NrW17qt6Do15L4X/bjF1LHZrvgZoi8qFhRY8hWfA91yhd
5dvZvfg0jygTNfHsligNAW1f3AGe/j4WBnZC4HlCHXOQTXIEL6/BN4yq7W7iOUxOkT06Pnon159l
KfzAo/E3020VdHPxB7pgNg3b7OK7PnBsGczv4ySuG0fkA8yyk9tkSUwUnbq/KGelgIb00yCJKml4
pY88ASYv+X3wsqde+3olZPoGjFJvmDIdYPv9brUcoigV6eD5k6H+mTKUdS4Cc58g6nAYwz18vp/D
a+vP1S+HjZJ92a+nKDhpMMcoFQl13hVHFdQGB8q7g5gACHWwvOixPkdNDEg3W5DedTFJgRNpjG/W
q8qBc8TEyekVhVN4aKHkv9eyjN8zYnJhitCiTtKeZpqxQ8W/hOCBJ0irZA9rsosxYGD8qsMjtL7b
j+ypOtgUAmmmY9Io+e2sYJhBJb2xlfJiLjnND11kExiXIlQnwydjOfmc0WqKnaAxqq+1t+CoudJN
HH/pB8PBYXAri0C1dmx3d11r1TyluMD8ZzIOW42zLPThJimYlPbXxkrQrROWpGqEV4HxySHZhiyX
NRRoncfT+NNa5FwAq2yXxGGJuD304p2Yq8SP5lHUFIxQ003qtisIpLEVv1Ju2awb/n3rq0IzFRE2
jvFguVlzMl8oPFH90iDiMMv1enLIPjWFUC78+BeTBtq+//5fTzqjros46GjjBoaxkJYhX7KpvTGA
WDgfwL5OZU+CUyk4TpC0yuIE7R1mOoSyIVnLo4ditKAGfgK06f3AcQlIx8F2cVPA2ipw1WS6+pqX
7uD1xIQaDf1VRGU0NNpGAqzaP4PRYdGhRpgS1u3UC28BBjA9WgmHxtUwhK4ZrcJ1eEfRu/m0p0Gh
KEZB6iLTmAbZ7ZbpiKj8Edh36wwh6aea6NO09F7lyCZgX8KsNDbCduoRMes5OOqXlc4PXxL58tKz
5pbaSJlyRQIilg5SxT6MdDCFeQNY9139E7ICmrIXq98YwoK/ejOthzyqv4/zydbpO40N3cOiAad/
kXMyklov1kaWBnGrSam4pftfbii2JMQ/4wm5oyOYyLXT6z5Kve1mKfdHARX5B4VXP71f3pH8O3B3
h+0I3MG1wYVi1UUqxi+9KHUHivaATQhuByz/iKgqtYh2CmZTqJc1dewRZDk4unTM+B7GDtX+fNXU
VcA4Z4tJIFVPPt9AhG3m905tlEv6ALhHoEzHu8FE9cjj+p7mAuQcv3NqwFtAjQeV6akGldv3Z6zT
MhFgYGGiE6G6pTCxfaBmAI9xLXddjzKj8yLCVZlJpt5a4L3iRtCzDaSK+n+8k8zY8lJQForJI/iR
wqqBIiJrxeimloEKzoKM+fP0HfGYEuhvgMkV1YV2pFqD6VaYctI+az4o/bzCsv/ds8SGkMc6BqE5
Mju6gvhqHKeZo2oOv3+qSDzHt45aLqoiRBdbMKfMBNd4j7BCJ00YUhh3wDxs6fJhIGL9ysHTPpnv
PTIVlVWtJEFLAIFkSHDx8KgtBbP5q+bUaZIQu3SOHYAu816zVcQLJ9nKcVkd8sKhVekXG4oa1xo+
Is9TewWbNjNjuCDNMNmCpHKTgsndPbSVpcSWm70zdHihJTux8JTzda2P16Gpr3W5GB6gwjeiOKtY
ECvS8lnjkWFaUbUwPLkitlI7+0APrsapy5BdMg/E9Kx+lKIk7fI9v7HG6gkZvs6l/yqVsi0P3YOW
bSjCLPhO3B9tbEJsq6L037E762+g8nxaJSacjJOPYrDLkZWJHpggvtqWr4I+0keDyVNVja5Nv4On
SRAuzy2o8eCZcmyaZTjgGz6uM4tA0yfKpIlYUgqNZ03V0j1WSbwkQjgFZn3ItBwTPSdrgMm/p8rj
+n8Seoogu319Rz5MjZNekGF9URs3d3ddysMMxFKF5YJrlf/5hdZKdVdQ6SuGzxDvgDFj0W/2TlwK
xVNX5MDSVrIPX89t/LPa+CEfnaj3SQcr/abyubHC2fO5W65q15jvEcVlW2UHhH2MXvtEJzaN7Yqu
YUw1AjFbiz2wdXXS+ZYUoa1SAnR1cHDd0nNNJcXNRazibQ7emF6j2pJex+wsNTDKDKj2FrsV53e5
dJIaNvH+2jw1wzMj67fgp8nJ0rrfgmuNHLwwv4CL+rdXpZuJOqfhHTTn7YEiwboO8BI3SaSvxi0M
rmxhfoa6450Z/TPvxYmX7XRnQAiKB00lw26L7x3R6GbdWP4y0bDcqWf+WVXQtabnM18eX2Q+MAN9
HZwL2o4y+lKeEXKfmcEONIvfztlYxwxsxX+uraxknOr0QpvaQh0rU7b1v5CASaPSqVR/UCvTcvQw
XwejQsl2vwZi2TbXch/TOlcGqBVdsTL3V9Yy5SoWN3P501YvfHE1VwvA40JwkdVw2q0kN7HbFjGA
zibtxbUNIAryNpvN8BXE8zxIidBDnq9MIhtn16V+lC1EDejegLy23IDeBd3I57HjUvaqg7l77Tjg
4wTTZMJ3Ld37301qpT33KkWBzbGaMu+i1nGFo96FdqEHDupqbeonWf1wtfmZE1RjaOC2Urs93Tdj
J2/pilRbL6hjtvz6JyjFuAKy/FnSpiBAENNoGGBYPRuYlSU0vxN/ST5yjozQqW+t0ga7bQaDcOqy
+NtUh2vLh1UU9h5CJyy7rMly3vkzWxRfjjcnNyqwe/VbIQPWyTANdIipRnVXMuxMU44CCzMVb7Wz
dwBtUwSKUjJQcKZ5FDUwIM4bUfFFTutSUUUXMgsArkokian8SQaSeQTrcq+tFiX5pZFtFa1wM8oR
t3ew5nx9+e2qXNnEck4rne08ikFOYgF2OgWVk8LPpKm1Q33Job2TT5FnF46voIReqVfeiqz42oND
MNS1vAabg3QEZBTMLQU7W2fxpUlcsnmZfRl7u1f3d+0niutf3HbyRKm759oDhmtyA5HcAgyonFiH
+jm/ou90otHKyv6RYmMx2EHy+h8F5Gln68QtE/J2GEdkTZgwH0I1YN671KrXN/jODDxPhM2Gs5jE
CJmDEMdMzYliyuznZ718/rlx7c2/SWxfxeXBVhyPukunPcMBm3jYW+soHz6QEr9Mm2w8kkzlYOgV
OEbtyVYxG3SiFi9sW4bMJi+7L7/pMkhlFmJPssYizi31zoNVd/4AV4AgQkvL2hrwmDfjQFzXU5wu
oej6Rpj0vSBjP+Sf9wq38vrXT2R06gN40J55ISLCGQFMVC+dqGwV9bolocaXaQDflnWqsAUZ3hf7
ya2GQgZ91XarzA/DcWuo6Czg3S/L/yYI241EAPZWb3OuoWL/JWEQ1X8IY3ZNOHnRnsL82xtxjd/T
3WOWwp7OLpgEdub3gFXohnSov41FAKMizGtrRErR6aSvNC0n5caTvxLsa1H2qtN7Uclb4XQw8CVv
W/zsXVtmi+Uw/lEkRaOLfCvaoBFClkPwhxgT27k7AtJ7I5xPjZtkd2Qoj4Oa+yKAgswgJG65I5Gj
gqn3uQkd3WuiSWz73AdylNsOkv0S92DYLU3/t6qSSVfuxJvzupjavqrA1ZLuB/i9e3XFz88gB4KP
pVweJe5UCDXOXZg8tCb9T/bLzngx7f+AL82cp4trXiOSMcNFeJZXD7hARm1mFS5+e1T7vncdDljZ
36xz6dLblKmhAdIfZmUtsj4s2UbjJyYyzf8LZ7EamVAKffr4Gxic8ZlU8+cPY92RFHSYlfdXcry4
pck8QOy/KnukDpGYeKPJJQKv17FKQ9EPNYkqSM3nZs6m2oiqhEMABJb7NNER9qQU5fDX5O+RxZAs
0bzBsjD5NvgXE+zTVGNnzhILEKgy1kx/mDKLruwIll4w79rzXbEWlg+3NA5k9bpFCIz4YjexFX1/
5HdTGLtM7qzamlhG2t8QZxu9mGF2+/JA0Fliq3Jn5Hzp26xVX8XPjLm8g7fL7NTTY6B/wwmUt60h
wTIpXOjW/esV3888g6lNWuiJ9mnCUh0YB1PCn2Z5Hdfv2OsFetI/265fpZRoVLs7iygc2+GegKUw
lL8xwlEkm03HiAEltka0eX0gXMy0SW+I4qZnfIvMN4xxjnng2BgZldRqEoI35KEnKpE5yuxyEVj5
LnkHe3vDYniuy3TiOoOKrniW2VG5dVonCHCNzisJEXiNg6o1ZEgsqlzM4eUkGeTkS0oGkdj3wP24
vsg2eIdOWIvXfoWn6wTup7+OJ71VzcOL6rVnz1MljwVub1U5JOxv8uaaktt3mRKw46fP43elHMy4
4BsI4+CS8AHYrlrUsQxl3eOb2tBBaoyFQ1C2Neg9kyvN6NkR6qy0ebD+mc9LkOyNgnGolzX64qaj
Z+yNBJPpW+mwiP0S/FqH9sIYRNnW44oL3HkjYllykMd/2AzLakt56UfLtXEj3GWn9EJ/anwWIvfl
TOY/P/K1ZQn1LaJcP6BsugxyPg52jqSSmO7LaN7wbj7droZV3C1ayPijK42RM9/bpLEF+zAj/vsn
3gm4Xchq0ymPv7W8/lQOXrQCvfNb0ZHQ1aDK+r2lnxd1E1Tnat2ldkz7oYaWHLuvXk4mVOsNsKyr
iUzEkqroz/5J4R6Y0eRl/Gft2tk5Rnlb5LKGBuJMesbXCx52srtiwPlAU3wJzq10GuHpXJZplsbl
JCgFQIWuF/VyMxC40Nw2A2ZZdn5UInqmBsSGXnCX9C6KvImOkLTrB4iNK5TZ6OEwsnycKqZxeLdn
gYqcDl6KoiePbn7Or8nLYZdXcRJmbDMOONwa7UaQycwoEHPqkhncmp4Ag3QG+1TP3x7s8VT2iKL0
Gs3MeJbpqI4DgOLK8fAt7IY61wRUk6WEbx1QuN3NBfewGkNpXy12xDF0oCpvMIurAaABpqbpC362
r5q4tLInj8YJCxbu5uyHTQ0bVmfmHc33sPqonrUBX8J5lCO693pO5rblLScM6e1Gzc+UO6GRZ7GT
zl8LPRL3Tu8z7+nUFlXTCT6aPM9pBbqaspfCFlDktJK1RAI+DPPDuH1TCc5Gwdtmgtve0POpMRht
CKTa1ocWICpVvyYQ8TTvWSfiGo7j4bLfvBG8ek6iPNmNqW8Aq0Pbrgw/U72giEIYieOUS7jsgQ6+
rfOq782LXr71UHoX4ZZFeZj89zi47BA03oQ6NRqz2+1xAnwMJXg+lKtxZWMAC7jnUlr3E5u76m7+
cxkUSYefy41ddN/5n7kbmunsgQLOkFxeQI0uBN2mZyn+6upt1id21YT6exKdVaWpXYhvab49IGyc
DIJPWNJGGMLyeF0BFjXluwJ2jcPlL846t4nqZJqjxm2zQoKwMPafd0jblqRgNjed3n0NZuoJyAvz
rLayoR7xr2fXQRlSnwwvviXFqUJles4bnF+fsQK9zBobsBEv+6G7RWBbrIV1cMfk6XhMY8/Ye1BD
31ojYH8MYiPWKqi04aIr5jJi/TqaZJoNdhg1IKmMOy3bH3vOxQyZstNUx74nUfVnY2OJFWtVCPjr
fxZmTBkqyi8VMn9q14yrSb/qFgbfV3xtZQfbeXAvwehzXIzudjfgvrEiBKwUvP4TYxRf1tkdwWV6
qmfHmpsmSK2CkFhlFhFBkf/9XDy5uB7rbZkZMVJ3Ou+Zpx4u1lqf6chrWr6mRMVwy5B3rqFzc63S
+qi38EPouI71zfzh95tZXkfYtISoypLiY7yraJczL5kIu6gcOcRhqmUdurDmudEVEpnDkUqyUGIN
tujj+2Yz1eHRWCI5vybQOEiHqBOMuqInjvLVuG8vcgkjaME5om1utvq8SXGPp+C2IXwYQIUOQZ5o
mtScabtPDoBOtKl3As1wb1t6KnnkMsDlvsFPRQNpBHinRL8zu4lP6nIkDPP830XLJbocGS9uiDn6
B4kKc/Kw0X/cyFLCCrVzRzvs/KqkG2/450zYxw6v1gckCeYXHcgEGiQbg+ELsDQ6mKoH6AS6Lab6
+783xC2hVXD13CL439Zb0hxWxWyRxw2kJHUu/9Wt0GWeM/gMzU1Rgozn7UooWBEXqelVgzuwkS0W
Lhv6sRwzCoFeIALLqNUvp3vPKHlVHz+zuedLY+TZxwXFq7AV0+1sybHUt8Jb6+ofTqvNk2kFnx4M
PE3srzsc1GQLKXlA1erVbkEY97DQoa/v60pCAqyaQJbdLE9b/IwLtcAWCyfa7bESqvE31kRRYj4r
K0piTPPD1Ndf1l0ccKgLNNPZOntimVQZ9dL3wlJCvJIozqqMtqtwHJgLJN8dBTcA5OzMd5HKOqK5
n4ams9Qe8yyXhb9yWHElOQzj8ScOVeheAB+uDv2Y58QhUh11FSSA+V98ASlbGfIZuozL/FwPwk4G
t6N4N9a7Gcv8MWxA8iEplt7YAO9emsCLtjeKLtNiLq5G23Yx4nEW9bw/rcqDKU8iPt03Dzqtzcjl
zcyVjCzL8cgx6vtF3qp6UtsggDpDJEti3hYk5lF+7gSB2Q8N2LNlS683Bgp/0aRIjI1LpuXSU+1r
bdUVs+QghD9VriMTe9rMRf21uwz5pTE3iVE3Johyg70E8bxxEgk3JCcHIPw8bj8ajWGSU2qYM1fr
PmBvlbdfLKyumGvTcGq5ewnxHbX/jcFfsbdFycYGMvNZt6Ek2nvESNVADZhbAKe5yGKaT/ydQC9e
liWOuI4X0aIhXuAYwT/q2WH+XVCYrX3tpBAwkG1lSMEzfvDdRfhyGtO3HTTS/XiOURXYZzMfofki
wHVzFNcPglCZof/whzOKg7OWGIhH4gz49BIkiQSIl2dNQBJ358vhi+3wPSYKDRa414ECZn/Ppke2
aABV2oPOtiS37t0qXqPTJSdiN21V7IQJ+GhhkR8kmE4/F2NitRG/7PWgvcF0Q0D5cM6XKkd0fykr
d4QneZqPgNWMLCKo3rA7ffzeZx+ETZOBh5mtmYKsQE/+X/wVsUOQpBNQmKLh2xAH7goyZwRyDRB5
m9or74bcisTcvpv6EFr44AODhVvzl4LnL9MuiEeOir2igRPyilrhfjmVfya4omk9Wf1yyI3AOEvs
gIDEJF9mZW0bGIzIqevmCDJLfZxDYcEKy8eBAA2e8pa/phL2uHAsbKZOGg7CU8SCcwYKNl9dRsLt
1H2LHnPyWNcxRuyBomLEw8WgP0pbvanzgTkobfszq3JhsZgax5OwhSSQDazwdzQD/Ug3mbC8Qmw/
527D3KVLcEYSHfUvaWx09ryP0y3xkB4nWdggCF3nKrSEyxcqDlwDBVSPoRrQnkEFBnCDiYA0565r
VcEetYR6TqBU8ipnhJnGem9JdJa3Uv21W/BgemF2vXKO3uvAjpLKsLI+g7eYmac+/P2WQJPiWmUm
+oeqi6p8RgqFCn+H/59H7dly1OBFnqOU0LAZ/uUoGDXvxEON4/fr56824D8fEjLyL1TSyFwKp050
PdKcCMMHZRvP6SG/B6KaqTPrDCL48OY1v6wLZtTuOCdAG2Zdg/dnMr+0GamPWesMiO5tUt8E0WgD
5JI0RUNZXsMPA4gSf7zH0vgG1FhOBcJbrWmCTywzIoklPvZasQS+zJRYz405QH97G+n2JQxWVwH/
YCwCLtxa8JGbO20XJ7eQHWNsa2H6Z+jDar6XMOEO3egv0QglCBTM2ImD4r9TZ2c3cAz0Wev5GitW
WIwt8YnXIUDhnsCQgsXqVNBMdmIYL05dzrDGdRDJm1/jJwEVyxTySWhWdohbKuC7Dt6yFMZz/12P
vLnSFxL6mtOqRhsSMX2mh+twe73LJEEdFQyAFnpnhL1MqRwxQoXi7uC6VQMnfIUdmFmz40vTn52f
jFv0ILSS4bP7l7Has7Q0TWm81ryKGUeLiAr6EskXiKKaaMy/JqzsJLJT/Q5T47lA1qIzqQ2eIcJd
abF0Q/9qRx0edAuY8N7qG7HZoa3yrhDi4wDvmrKvMNeegdg2WJV5BWOwVw+vik1mubTeod6DPr/9
tQv4Ufh3g6fTANiC9E+uRIeD5uglfXO9RD4+NSO5CIEOWNwI3ttgjIsB4ncPJHpH8TIS1Zt8Kl+H
/ayl6HUIlmS39ZNlFOPxUrNpKyt2YrvjUtYKQKAgcAPnGzi8sVMC96bOFG6T9ISUxiu0zTlRfbN+
9fNaPDLnKKoneYRJ6VT9FCae+8nacVkCbV0v5mXUT/JRFAcdp8KPGMGni4wWBrXKCQ4uw+nsM5qw
4wUzKsLgt60YLj59rJabNdDbKzRO4YRnB0jirsLVZEfdom8oq5oxG28MfWxj3N9AJXd6Y+AnrSCu
bOyM3EZNkDbtHvZ2saRlLgiXN+YEW73yKE4b+wmavsqZFF/7B0PzS5xctVrCWLWp4laxerimgn/d
88K5JVRGbWQdLPmW0/BZ/BgNi5hXmMdUsdEsQ739Tc5togJLD442pE3Y1PrSZlq4lQSwkiX5RkCJ
dYqLDLWH9NAvOO0qCdWX0Ck5HnfKEZ+6U7TXo+zDVAJl5rzrlNLeEPgQgwlsiUqxJH37ih89LM6S
MV41hp3T5eajW6DZgeqSC5scNajNtTjcCQJIIpv+6PHY5cH9OnM1hJGnQIwr1qlSVxLPms8PSmDq
FuD7AXFYOHd9CGzJ7awz9m/EQsQ/jRKtpbxILTm4vuPHrlcTr2b6xDfe5KudjANp19jpmZZdb7qY
ofx/3BFAbjJ+T8fZoL2z3HIcOAVIZBHbeiOPHqvwoOfnTD0puUG97AFY9cAQIW6r9SHeHjiX3lmJ
VtM7Uy4bfuLYFocIrBqGo6uKGRwWNdr7zb3CFQcYGLr0nH9kXe5wRZifxu5FYZFaE4cnObo7i1Hd
pTBPX8g1iGvlbgv5JrTTCJB4AV5SJNrEZxL2uVSXUlDbTXo98j+yl/zvFdjBJ8SVGwcmffx3XE0t
LdTkDbcwWtTF/gNedgyDe2NMuJw9EwhmTlISQEhXkzCPXFkiIgW6lm3XztzQOQWPTLbxcuN9kRDp
D4bbABwj36sYpdUVt4XmSv3LN3PZvgCPj37dFo01jPX+8vYcDm5UQoIC2VAPoFtnYyVF2mn0Yg6u
zwkKdPjvOn/Ysl143k00F7U7hKH8n0xATsUC45TY45cTGBDUn9Xtj4JoBO4xmrLvLC5Rn3/gAWp/
tShMAqRDmtSJG50pj9zKwOQ8g0QEbx2YoP5Ms+jlhQg7I8ShYXyEsP8qMHx315yS/Leg9GhZdmwk
sGSwTU7AdGhqLO3fI4m8ZOPS8tqcZXo7y30jJuu1U/e33NJSDIiMQQpJ8ON51zHb5taNn7M96UPV
Xf7l3yBzeks40o5PZuo7K9Ua/Fe4Zs9LDJhsptLQWLzaMms+W+ZWGsz6UBEAbXTOhJooeVschLQZ
nEYHV0dNziskKr6zYtHdz26wuZQisSUNzNbGORzMB4FsXZs+rlIJcT9M8vhIZcKt+J6HUpNFFCyA
2WfnhrveTEF5dhMGuFC0dxwfUsiJayW142lrcYNly+6hyiFlelFdLwg65QqEDk9rwUgIeXaEIGTM
JoW2yOXtZtTDYMTKDK2b8PpNpQ61qRLWlnnoP8kdJTXQILFNgQkLmtyjlRDMMgQ8uGKrGKvBgHdc
Cs9jDXjI5ErPLuMo6s2Pga59gi9eJFZ7+NkLl0DWVmIqejMHMQrSGPBaWoER7zt6UX6TURzEF+Yn
NNvn8KsUIqmmhHnUi8iO9DNuuKVxfn2tzdRhqC/rURckTRH+fIy6bqnC9orVeIArNrY9BzzGWl3G
PGURjiiIHK6R57XoicquhuY48cEArolbOLp018+CErqJk0IBbH0PPPlBnXb/OQgjwD5LzhAPiIfh
VFIKXuwiVio/h7c9TKwIjweKWv+tfpU1uTyONXgfO2zwqBddG8euYVGa0mWl2rVum66ZMogb04Wd
6dYvYbCmNKvywRPcaB8AWabME8DE5+nF4jdaK9TlcsUvFbsqwuH9QWlXr+/teBhO00+7bzCbiaN4
j6xv+nTqlfoc4/tBBm9SNxgYjAQFqmlr4USXJS9zbbLup61hmCLdKag3LWL/+jwtR6LBUfwhJcgJ
ykGMdVSZjaECZAMBjGjRCQV+6fPEkr8q0MhmhbPoFFTkZ2mkwkn1gWp8YhOWkLBREcOm7uAiyCMT
Zcqr6vYjxz3zY3Di8o/HTMW8k2J+SlrX9o5lvHsRVFDKLqXhS12ZCAh7kMLrrfh4LqCgAaNTELb3
njywMpLSCKcV361K7wXYWyvWqwSyEMgV8ljKBWsYd3X4XT/QQY+zrSq4MoTj9oDMg23H0iu6MUUu
NHglm5MRRLtDqHMSkiEFTgkzA2ZAKDDj5/ZIRDbfHYro0WE+eMb3U85V20lIStBgfkg2ZBpnAfVU
25py0UD92vGMxQ27QJGEPbuEmpXfAlGlJfvMoDZehx3krFdi0qQB9JgNiZ/+j4xMWSoYBQHw+ak/
gH9bo1FyWsThbWPoOmYqEevgCQvWlDKRJVqoW4JDq3JYbSAqtOi73hZ1P+0nV1Si/19mm5o3hznG
E5/VOKFRbFCueUtlvToOXVzO2KCEba8yJoDnKjD5bPGx7wNmAelKIUsGIy5SsEIVZnvfrMbfEeTx
P9QqdOTrh1VOkZ8KDRZS19FhuWvjHtZUuCxEUm8mC4/JD3iCEENtHR/ZV8bZCVRLKG9sDN93hkl/
ARtSsB9M6cqRjST0WflInhkqbyMXvV5ziCiJ2V4uAcpUIdINXdMuYSOXDNcB5SHMUF6LXWicfq7A
cNZw4bHOKtGU8SFGHLC5zDh8BnUefrNOZ2xKXJ9JwKiwGXsRjwKAY8UrZad27N+TvJFmP6kqtk7t
GNEbKH22vq2kENi6bnKCfwehxvkpG8eBfQ0JpdNWBirNjdN/dKKcTYhbuYm61x4fafaJYW1ElpGe
QmCjmpLojrQ4INvIdXXwXTiTYsmnzUrou9A4OuTvbgXNo75EELX1LF8BQFLEmJLnl41fR8GT8Pvu
LpKaSX/GLJmjKLKeaP+k2VZaAgUOOx+YUMtLY4ASJSdW3+Dsi6uaHca8Hhklj3KyxEQyhqWeL9k7
HMhs+ZD/rYdjpWcDGSZeHNej3MMxqSDdVgHoXhVuznHyjTOHnENrOteR63Dy+A47ph8aU0dt6xgR
PitnXBLUtNJVphgY0nYcOrkWOSZx6Sg96JFFUPfUDeDD/Qa4gVGfBRmeBFiV6R5XsvUgOrRPZ/Qw
TKOVVrQQhwCG14m3MFZTdQMFZR5tTiGfIq9bGT5jKZGXShvj8g9/H87tt20NrP2yztAYKjvABWXx
eu9aZd079XA5l5wp8iS+ynSF5RlUXncKwI1TmcaGbzkFyz/BMuGe47nadlYSdA8y2GtDC3NQZFu3
4kRw13UfB6m4UUhg3xhR/4zPSKBBEyzXsECjK20/PywNfDdulvNBWfNrA2uT4R3CaWrFTzm97uvF
FMPN4v3uyIcVSm4D5hivMFX4i8fU0YmmPl08Th2iCXeH/kqfzPIjqcHPVvzyavN23gUQreWM5ArZ
nGV18+yfwBFeHi3hwduFZ/VsvHKtAiW6Ko4sD/o9Rm1oX9Z+EY1wGeYOSK5MXrEQW7OZXLCc6JaA
LYi9mR01Z3VkhVkp6eacy0fgAye3mu1nlil0uRlTa9AK8gR9BFIj8U1EeSStkF+RrcDBrxZn8TJ1
ZoMqrJNCWv84RlTv8MIO39uwf7fCkJSwzY6/A3R6rEzC5L7qtMzm+J9TjP9d0itd/tOXTXbbWO9o
050P+MV7l0IJIkH1HBac7Jq2NP/HL+VPQdkbSLSZhfgQlQYudod9HKFdCJXt030dYVKf57SjyF9I
9k+TiE8ZK+h/sfnh9g3S6/k2nywlw9LdJ8dnRMULB51/6wBNp7WsB85YTiBw2w/IPI6EtHlegWIj
K87xxBU8X9g9HjPykWrX80CoNP3u+ZfGzDkQP/6Dr8UpERu5+rslL38XrweHCgS1H87WCvOHRq7k
jpP4S9pFofwvRipoMH9wNo4UBKZhOPcOqsfwwAS1dQ1yABUd1TFFKbDqS4fUCJx+d7781jXO5UBQ
EgyGxjdc2wz57CDzVo07DgZ1BneoTwydzh2ng4N5ebv6Uh5ekht3j8/6zX4xtLhFM1NmncJugLo+
NRBl/Emi5R+DbJ+0g59vUi7cmvBWUBl4TKq3O2KLNadBNnHaOIhi3tJLRwprDnoD0r6OwZ1ATCkz
AyE/w7xlFBMEsTPXlDJIFTBzmn9UYH2e7fJiv1frkIs7qIlU/NpQNHUsf+e+W58+URCwFuZZ4DYA
n/OnFcrRs6LrUnGjlEX9Y8SIV1nLOqHp/3r6/eQMReolE8iaw4mQBxZb+ccTr1bkcI58O0LnKWCW
kBUzz6q1fBsTEeR2N38hOEHOjZ4jyvPQXcLg41ygXVHsuctn4OQ0w4mwIVe4GjRip33UywoD4Yqc
Ppf16ru0vdZ+V0PDcKDH6T/1srapVp3UKO9F8Bq5UKqZBULDfNaUd1DHTMJmT2/06XqlR5cTzEAK
nDVogaDoR25ql9EXViLDi7x9M/AkhniaZdPkO2sSkzFUPyTlv95m5f6QmJLnMT/VLDiYE6X/Sorv
+xJ3Pc3mMM++FJq5Rxgd4HaP6PeYxE/FAV/9a8S6Ie/Ic82aAd9fA/QVaVxk74RYs0GtPqz0f3Km
gZneE3rPgON7ubU1foo6zSJZG6Y5c4fxTuCmoyQIxZOFHWILz3mWfnNNh/imR2rn0eQaOKPI6i5F
hiqb/fAkq2i0oT4ZpBbnbwbvws9WUhUJe00zcBZLGPzoJBmk0K7eiAt2JdOcUUpaYuXSHuhQg2XB
gaVd5hDZlVsYLtodrmyIG4+G+kQCrMsCoZPXTxa4OjUieXUIutXsdV/dNQ6RJ4aJ51EnrKsi99BF
kBhF5xufUV4VCYnup2n27jAeM/7hbo1Qx1tbcpS38t70XgnLsEya3HFSZWOiDnQLjNeThz0uMjkY
Lq+SjYawU7m8CYuCUWERgUBKM7sN8wQ9cQlM2sDN2Zfx11ZJ+h0zgxXqhQ1XFzyTSCaf8MVrBbvC
OKH34b7khvw+FMbUg0n/O1972VhAV6Mk0MIY/WlGOmV7ObOhihQidjFygz4mB2wS4QTXn3z764pr
9OJyFjovcRZ5k+takmCzo7LidzvpFvrYpD7gFZ3eYKyxLwkZiwDgiwIT0WIX66+GZOyiPwc1yrRR
b+gVx2BLaxcZVdDLcgvVkTwESyGP48StETA4HqCsYu61N68frFdWjroBujj681Pwat4Y7oK4DPd/
rJU6CulRyQnYOlGIiXhnBSCbIp1BhiQWN9ZkTF9KedByMKg3rVX1qKccNmtARg6eATDWW4WV3oyb
CNBRjcDCw9blou4IxW3lnC14ZQ3vy7hky+echf5ikHAQlRstbS6SDXWv1ji0S8WORMuOmjPR/xfF
WTTCaxc8hGTUuSlmAxHCHNsYbIpvCVqmkxxQeXMH5hvzoPFivTm1N9Wvn0DxR1bJSABoElKZ4wOQ
AFQavB70xmaHBe3cTRBId77xR905ON5Px+cVDiFshoyNQXK0CdgCBXJ+f57ygHxcNu1+w2iWXacv
ZkYKRaTZ3acu9ni8vqXEP0ZHDRjhsNWzNyWzs/rn4dBB15Lp7cHFX/HGnDEF+HH4gLVF0xDfmC85
F2CGV5ZQ8KDvp18tAq14cEoEbgE0tQ1Z3P9kuBbZn2U5NmKSuXxLAfmm7H0929SoVpqAxrr5tFFx
F0xhy/r2NYd7ef0mT5tqRvOPOCLpVp6S6uYZR4Eyp/9zGaP4P1Ez6JuuIsG3kF05tMHBfsk7dGye
SGeLDQf9wQZduMzN66xhBRUbPsogn6cYVVf0rR6J/tQ6Hfk7tzkn/4pZfil4sTmsta6gsViwqyNw
VhtL9FtTqtdEz9DMaoI0/XUkX6N3/zrA0vrjX02vHTQVtW3W6wFSe3hViq+1BJTGBePiYRALUPi9
XZoCZHkjuOqRjhOTRCZNgGzWZfNrLxs0JFbiGjTnzRdZNLdysMV1+E323Wy84OAmTB2YPlGy61s3
lUh2FLLRfJkL5pQllwKT0J1BqtbKcQc5a3DW7F9ljrl7wOvH3hKPegA9tOMsFJWtP9CyIrlNPrMd
PCVdEud0ZknmnAkk4UpwR4H9JryrdVUOZ+tN26n1gSaWLBYwbyXm0VbkCeHIRU/NtbVKBBx0Bb51
JQ3RRDRd+m/3VwimQYA1tmu5b++rYI+XS8Cy6tU25VHm2iERy6zS9YDIl2xLmsupRw9rRS7pirqn
UiZAskhraGqeMJzy4XLMKpRP6FmFmvKWzknkYcBJc9JiNsbSnCBdP/QWGlLFu6lPf7n/oWgvm1cG
WaAztNBdnAJGzDDuesCstPqEChBq7tD5837woX4rb+lmr9e0I3D1Uph43G7V3R4OH9q3oPMhV4RV
mTL3OYSlYnFMNbaAXl833u9auV8I0GHwxCEvXytRDFaTtWYRIraasPQvQ0J4WJ9S5On29uu8V+XO
xG2lPScVHJGykj2yrV4QnHWvkgMpY1VNDP4e2HtyokQ5BYKUWXAIvG9FmvP300Q4MOasyezvDhI5
WoGTESv3GbX8MOjNqO7eWYokEF3CT+e88hQCWRvnh8ZEiZcIhImx1sSz7G4jfn7e2D8LpMYwVWUI
GORNsKMl8FoVROmeNbe4emDyjL6BuP9T8OfWnmWXnums3D3hGk7ZYq9MzUsxGtjKoEvWeC8ZClpD
o/wt3SfnlTlCDEOmG8bl69VXbRA7vuGy5GeYjnV3FHxpiJPEgQv93qy3EqP1ug03nUn9Ipw9L1IX
Jnl0zNLeufHt/jnvdPT7TLiywWQtoOit/XQDJyjUx4ZvTNuYnNhm4wjrpUuxlLg09nE9y0Ueql6i
DrfMe2x7M4ZFGEuUMrinVAPkUIlylFbkPnHJ2CXvtu1XW4Xt7e7VDri2c/LYv4LxRNOCh8j/PshI
w0bTLhAkXGWzDOCJtvjx/OWmf4g3gLr20B1BhyD6NYdTKYU1vik+amg1tv2ddqWvQIldrb2SpiRF
HfIutUfKR6SoGWcMCWSisXh0XpP5HxGU7+O2mTtaT2iSpYINZ5hfvzk9kC8zqglqxyol9nlpv+62
vrQfcgT7JE8yoWHHcXktwYX3LsBPQSJ2MQR/koPY1ux6D8vAS1cNwz20FTwjwcsCzyuRjI/qi7xw
akHqrdILndOY6Zel27G2mCEzhW/ZV7wOJtlewcTsu03cfVAzgYliuXUfWWnz7faDSBLO80UQLd0f
a+IcsWUWqKbsXT34RLZ/N0mq8F3IpVA/rM+nGcNnIh4VCdYYvLQV84rk7A0aAtRFh1OoDoU52bVY
4f+sW8xO+BLsh1XWcKClBr/qgOETBG/+Oaj6MFhudsbZ+fVLhMWlUxQzhAJJun54B1cmIMr1AXro
BAvHj0yn/5iVx8QWAqa+7Rorhcj+NBQml17CetqTar41lZuQcWyVW5rSW5uNWLYvyEopdhi4LFjW
6UFkHd+O9ouRv5DYzbc9CTL82aOomfm/9t99S0w1LXODHcBtlyulzrn1VF6+8S2kWidaQUU0zLlc
Y5wWt90OpURbrBN9+09aC2mYTRciyl/ogXkGNU01U/3Ref7XR7PgIb9STD8DdjFbsaICw3j7BMNn
tLocNGzNN8M/WpiBsp2D7HCrUZaYSvvJLPV7LQGJe4sDKn8DtIpP14XQOewVGH567yyl+KksC/E6
V3LH8GN4zr42/FWz9i6lGc7UbSagf6zXKVI0buhDDrwus4IxzC43LWzX0lg728hTyhUQ7E5PocZz
B9Z0Tmzj1K8413sdCn2FTDqPFE9siDhbQlu6XG4vBZCIB+ARVg8hDO1OePZnnEi8Olj47zEnYFAQ
6/tJk27QL7BZRpPQic/ouOGh6w6TNslqqg6veWQlria8gYsp3zczzvFlAFm5AoSq+HtdC9VPZkIz
MfhZxL6pyPwl9ab8CFb+l6zl16gPqMq8r44kqNigCLp5iY9OZd7oxZUBAJK9Ljt+vpFF0YXy2O5G
aStF/77SAXJ0T6ca+useawTccmjnuBByv9ZAcPsRRClZ46gW1iq/l+U6EW60iyLpuC6M8g2xp8Nw
IKn4WotvAlCmEwVf1Vqnx0zYiVVY/edtxvh+R56sJpRxFyN0jfLzViFhEV0uwGtHcyvqqi7g7PF4
nG9lyZRnLkcSGOyGGmIo1/VrhXmR2uIPM4dA1zBiAxV+3RnNETsW94x3gBCB0KUowJfhxHqfsiuo
n1R9NukqJIeaFs+mb/c9T8TNDVfETvvwN/YXgLvBGJw+FqnA2p0aRg8SLP4QFodVkNoezsjEFgG7
4G4LXtBdG5IZS5BMdpnUfgpeof5p+NwEbk2YZiRJNQq9X4MH9uaLL1p24jZSmaleZgv1XfmD5xOk
NPR0xPCjqCIu4WiLXpRPBFY44BNlgiC9xgLYIgenHqWlfY7UTiMRhNYtrwb1K0ysjS9K5KbZtovZ
T1vFQqSkK/30r9Iw0KlIpOjaFVXMIstQPiAsFa+U7CtKnQtY6MLHLDsZTmGK6Vu9PU6C+1qY+loT
4sQh7u/WONYxhUd8VyaBvC962m9w3qdjNCAZsPVMi9/ndTpOBkfgSs3AyyuMEfJN4aUzhJWpb8zc
ezxLrNlqgg4O2Jzgtt0Xwk5fAal7rx0l+J18pY77Wpp6hfwDpsfZ9zvfw7uZIqE1TXZd2jMzP2Fr
R3910RVRAvV+SoCyNy91X3ebqork8qPA0skZAVcfubsovecIxodZPl6zHCCh3Zipit9UpRVIaznv
+hqZuOUfjoaW75g239BHkbMmPSvSr6x4FNLKdNLokka4pIDD1oE1O55GzrLEcBAxXbF8XdiART48
zvHrRXMYVlqDrqi9MIbUtzPHxhQ2+2ePUY5NaXojyg/WZ0c3Rn3tjF6fsgOvSSXctkwOiTogyMnm
L488U9zS7qqV+P8EHUg60S807TxUVphlnP1yPSzpz1gmrKX/5e74xbnDi05ylyIt+boycR7T3YYn
AmPH9zyzVoHJArPJW6iL8ixZnEpGRWfxgaljLzO0ttzW7RFVzqgr1BtVahr3JEcd7mzD4JoJLChA
zuozFAK4v9kjvtJSRMwHU71mJ1olRs1z5QuD4hu8kLvS4srjv61/w8WoTDJWs6nun6ZTd5IeV4wX
CHtG6sOEIlEWAwPVsqSZQEg1tpgbGblDfq1lpJxQycc2JTDtGiLdJ7/77kHppFfU0/nrXVJfiXZ9
bZ/DD3LulMvEI4R9E0biGEiaRHY4Tt+afpODWl4Vs9n3fg0oer2WRQVgAUMMLmMg/cMPCUDwaqAR
oIK8zD2OciZPTXi4aoQVh9ptprwzhPEM0TjaEaEvlmfW+kMcsGeXoONTVCAOERmlSoAxrVo9Rxbx
9l2mENBu/DKwf16eKSFumMxD8lnZjYtfcyY+X0a+w32r4dgJ0gsCi+I9G3rclLS3AkHPWryXCzbd
NpzCfCmeVRtEC2xYgWnqlYuqmI7S8zJOKf6Aw0f7S+KozpyeJVV3/vOStenMKqjTL4PgeCh7c5du
aRTI5vIoSwd76Z4jkTcY7C9uwR0lHkYnH6f0Kr+LSn5vclhEz0WJO7f1c0k+ykuywE0BDbzeCMsZ
EEIfCLn6H6Ct3tvEyCWfKse5jDUAXoizGelj1eLYxoVqByzxNOmLnz6nI3USFzma0huFcXN2MyqO
eKWVwTdFZJwiStX/gkMkjW7lxsLTOEFbMHguv0KabaRDA+l4vNdIVQh9YG4EUJBe5XMfTzPmiSBc
FQSG8iw1ZpKCPmR6dyd9xK1+Ru1kibaaxf6UCCl767RFBFUFQnim5EpBH1lrqXZmLzuhDKh6Dhtb
oLHeV1z1jYfWIpeMNzsCrGvD4s0FcwO+xG7U0yFc/BU9FpPcZ73xri176kdLqNAwqC+0wCyr9Y2E
FiN4euIhEYTKSwUBQw/k7UghueUGUlwiDkZsfd/lSDJrAverzhCJIcbQ3vWGlU9klV2hC8EJ4k02
D1eWxGVxUB++XhUhutlUSS/hw6amGoLVCWbGPSmS9Gu+xJ+iQVqZSUhDsZ3LSCDe/7nTlCIq9t5R
JB1gN8B8gWQM0z8KHY7F5KW6GFF6X9DAZ3I8FmqjzH+OSsKrWNnzwc7pMAoH+zTQgn3wTvp77yP3
JU91bQs+M5HAaeycqNT1lEBYFCcf/pb5G5WeHUAx/BfEnrvMtNe/nxVjp9p3i/DPjTgx0X9TSHZk
5zKa5DY8trw3Id0YBBGI3g+EIC7zuzQqDMnMcudXP18EPQ8c5i0PhSbSULFozVaW3iO7jvr+u6fz
rOkGuScVOn9TXDIC5WukUi/q7ivlVlvILoTK+N1931DtLcXQkdwq1Ok7wCjDaY6KUIGh+JabAR9h
/hZUZZPWcjuEp7tI1ZA1SFLm7PN/yKLumQGLProRwl75NfZ8bf4v+UvMIqxmTHKxctYv+gNBm7uq
zFeVdurFP65FTZ9VeXVSXohzIBrPnOlkx3LIS1jaHcgusaeynTR4TkIrV+ZUxUVHLRz/QkokAOvK
z7PA2BaKZFjmWtCobbMtigmwXT4Wb19TZsXW0WXKAkM9p0zX0bdzsGPkW/jSPmEwMElwhOck5knB
GS6oUrxU1aP8tW4fBPE2ddHqCDEiJ0dOlrBeV+HHd8Gh90RmEv+i6jbVVEHtRF2mSxdweQ3PiBFW
tmCP+0gk/rj9WwVrf0ioamTEAhLVXvpr1jlhLkailgFpxzy9Zy4AgKFmZ6zRAzZHxv1rvRmf1/b7
JTjxKxwC9oCi36VbVm4P4NwJ0wV82XFoM4XCHItbt1Aw4LRD2EQ9Bp2hlbAlRkmnZqCs4QbsG1YH
w2plodPlRYeJyddpTKI6rIdT9xj6RyZ7qUsomezoj834MDPFse0kD6iZsXCQdNfSrdQkR+4RmL78
Xls1G8cluSmi83mmttNhxkGmKLQO7lOScHqj5RArJlHt1CsBuLBXqQQcxoW7+hny13nMUPYJ9J1B
RnQZGZGRJJyOnfgRKAWkXJT3yWCPQ6wz0pjvvxz+qXrxQPxO6sqCJz03DWrFiEAERJ4fRd43CPop
Q/0mizWGkS2nTqGQTH37wL48M3RorjRe1dVyum79Imowq2JmkWc6iDBAVndl3cnWe1EVzn7UVp5X
iQ/a6nhBlsdI5Aoevu95+eT9gve3Ixo/CctJHm1wKbur1gd6+jJ5A3QRMA3zrPB1wMnKiIc8P7s4
UA9g4JCuRxnHXp5grPPemRJhX3QZAWOgPCX4h5cM2Kg0VIx1wPWAmgJaSRMz7QlEiep5WfrqrJKs
9SiGATiYP7Maps/MAaE5DM9QYiE+IzIo2ARkQAK9oms0yut203DAODlSH4xNqJXsiZwKsXguPg+j
6D6llD49y/K8NA879QdpRl5GPbgXbdHNUoTvHEJ2ibmUZfQnrELsDPCMYaShdKVJvicYQe3rdsBU
G0wH4e4GRLsl3dqtipneEUDTro+VtyjgG0gvlKGgOPwKMjbxpDH5aV9kYDqlVqW/ZK8uZtnTGfG6
T93KXd0SNfRTsu4l5o4PVcf7K/aTiXLOezfDBaSx257cuZhay/QHiM5hT+onOWyVLGbcbP3U/EB+
bok0OWH1buo4+KeoUKHCVt6AcX2lXRyerfvfbvNYFTQLm4VcFN+VQ3LOYyYfo2dX8mxOh17BVmKm
dWHCitjLpzVFKWwWwU3NtHpeAFSSCu2DfUv9KK3IjQl89nV1TbOUoxsXa5JzGFwyC5/Xkv25uBwS
sHcZEpVDUcf1W2V7w7fv+OI5dv9Gd28zMEnBndpipEynH8ewX6WtqRnAtKEaFs2E36TBAmQ8gG6y
qmuE3Nwnea238I+wkLWrGAFNyAPk38g7BEgb28/U3CiDRKKcSBs2g0hD59Yei+8Zhv24JR+4xGD9
FKp5B4q5FQ3ft0LInOmnxCUnszDz++cTV9eloMM7umi1V+eE5f1jKoNeJapYVpEEdKE33GCjWF2d
AMHwPLUkom6XF6XFcFNsOmn6qZcfn0PssARHesxAv3h11FDHxfZPQNuB88LnyGrZY/qw+Dl2gUSr
kxswCD37mj4EyDSLl8th9WvDVZFDbzvv7e2SMqs2pWdZbA3h5Oml6gawm1jEtzXunGKZAnP6jHqn
2/3OISVXw8LEMsHfQLODubCZs3CoitDHTg6iSIKpeX7sE1zf3IdwqHveYAyZvhiyfjUnZ3LgCAe3
kPCWAd1Eu7pWLqziCKUx42Ok1Kt5Tj9bYK8BdWPsnkxQribEwYnc7SwqN0ujS8aboMK8kBDkSJu3
qEE33EvjmeLnALp451hoZ3w/upc6dnjWe1JEFIPm/shqBQQS5djLWppyA7epStUHIvJSrxGJjeZ9
+mi9E/EfCwsCnD/sgw0KaRjdppydicEg7y9py/OaP71WGseUJbHNXd0t6lOk8SngDZgEOpbWWFnF
qu78m7jk1dRtjEm3lUt7bKwTaLn5id8Y1PgDfmC/U6c07QI+C+BFh5yGGsQc30zJC3CLeC2RCOPF
sIvgpG0cI0TAkXd+LOP6PwLHI4hPNCne/OIeUFUA9/BbKmUQZVIU7cBvzsR+FWtfmqmyfM2racBY
kb1aHG2vEGFrIxn2WClMyMAngrbUMlS/12EmBt+2E5uyVpa2AdP2z96fSOPspaCHneC46DaNXwFv
N28NVweVMqchY5Z+mXeQpnHaTuYgswZFPa5WNC2plpUQpuHFCZNQNiR33eUIYkQ7VRp9i3EJXWLD
b2sXu7D+4iZCmr2k4juW+Wvp3o0FkRqGzLVqlIYU5FLvsqRF1LAm3ZlJBrl7qKz1S643rnkLfQwS
QaoVqto3xS18AiAmVw/EPM9EeJQFenQm/GIbrY5Y9IuYXsUxfFCShAqdUkijGh8f2HpAHFli0UQI
edB85zxAV6uQmPrtFIbmqzWzl0lvt3+NKnEtTNI5DfKJzSYrrJByFaZKSQLCpn6/sM+rpyvzjdli
T5FRvTaku3JfJoevthBS2eNfMlhIgLW0jr6uGemM8eboR6hZa029RuSrP6vrwDLz/dWENHSTMzTg
zu7dcFjZhJ3++GQSyYjohDulBKH+yeX7fETrDS6/7Ej4l4mTY3AwSU+ADuGouPEj3DTpMd0cy46z
pODBW8P95cdurSy5TNQ/dgi2V01cQQUC/96FWhC38JSy+Cgqn/hk+7q6wDd7/lXzSt0Jp1hw5HDm
BCb7GsurQEeqHPo8J6sOtVttxSyg+vtpmZPgLeXElpDO33zwDbGporWDH56jB0kgdJmtQUy7h0xW
uUnX+EvK82XJPeqQWTaC6a6sKUezcBqyqyH5S+4pHio6v9EWL7cQJ0oA5wS/81uSHL4WrkOr0Uxl
RmIgZWq0fS1SLa10Z5vNl+mJZN3nMU7qwtH7TGQuzAer1SdM7/F4e0R+Z3O62kjGBGrXuxatsnss
US+b/yoZBQkfeh/eO/9iFTy4uP8X970EFjUbHayE09cY1PqQ/KJ7wRb7nLKepxS21p/swh37xZeW
Hx84m0lS9uEBD0GSvwaMawa5xgNH00HkREpXC4xGxTEo/7JMWFavaY6rZV9nWRz5hU7cMm2vKgKD
CUYDXB3vNoafxtDtbx6OcPByybX2YKNL+lwrdDN5QvRQvOwX/tIKvyL9xlccILYP4euBnUetRoDL
2C+z71PuSwT6HIYVO69lIDoWpjXpcqCfBmsB1qM5L603s95eXvOoL2UnvodgJxMRY3tQWqW77eP+
IfhEyR0Lxtq3dFi0DnaSgtGMT5MunVQVtBzIYOkvLEOcIXcD9Tx35vwMcROkP2xk24C5J2ASB+7w
PEIVcak7bLA1N+blvORujsXYEAJ7oL11wKGFmIYuumGIob19pOde+2v8PEt+HMtF8N7/lUb+dCW6
3w765TXJ7nuP0ImD/VHJONFlOEdo9O2Lxc+W0IdPa6TD3lrbvj2olqiCXB7+SXLmjCXJYeiDTrj3
gdS4o7TOMamOw4OJ1yudlvW4vnzZJ3LYkaFSsyNBdZcbwWXpLj6wOXsdXZEPNG5SLH0Zv9eZqhDT
/LW5f/52KHjAvAr7mh/XDfbhLL6mNb8XmHIQGUAgJV+5kDUhA/s9OMyVG73GpTasr/xqsT5uC/GM
jX1CjlkufbEiTEgW87fc1jsGtd4hmICVjlVL1jC6maamA0PKzmPtyAHgcbQu8ShGMEsgizrq7Iuz
J26pGJgXlWK/q+g9pBWhze+ENf9ANnKntUrLsfxLmhd5BtGLX7pzLB+iQsjopa0rotjv8Bkm1OQn
ht2ltAcbEPlOQft5x+5gl5NXcZqIgJxeR//11BgeItkLcs9EMmVDOwvTJ+bsU9EcDSVWR6EtdYrL
9/JdccVjXTFmfB1jBJ2bMyZBbWYfaNbvQSmFeqp0dk6PsbLEa1ftB6NWBdplSY8nzLOG3I5zdZ2a
6Iz3BV2pIup//pzQfTpTjLSz9Ma4Mei+kGxG9mp4UiP1qLAqA6sdVSs7w8BYSCpO1g7oPy+G67U9
iHgQ0hjHpGrL+62N4U/SQZYjUE6Pa7t2edwDoMwLQ94SrWUAAjxIW8wX7atzPIR3TsiX5imEHiZ4
+feQZTD05Li2SIu7+/bvY4BpMQOe+z4JW8oW8LLIvISd2HSlKyLnqML+CjiZab0bSwi6vwjPUdaq
pjM7HhbWPUB+xESAdLPB7TO/fo5ArdatEHWipkccpLEJFAt/DMZ440uytOs6GlfP3Dnm7ZHzqGpV
2Pu5ss7fBfNxK0r5mdqzMrtMECCIAkLNdhzXdt3iaC2HmRKSYT+GnoTwgzDufOILdY+yO3kCbhcX
DWoEN5T03ZR7k7jht/n0U+gVeb7UIWJvtywl8tXUSkJIsYJ2htpHg/AAfp+L4NllUFiHdLtRbPR/
rnOACXYF2TlQCy7Y7+T5PfrdB0EnUCXKMc6A+jRhX1QutKqUlJJ/C6TiCHWWqPWjwff1Jyv1ATf9
B51hvDbzHdYJlelFkIpTXvLzaoP5+2XszVaTL/SIrRztvaXJFReXLcirxTyswV5hEbK3+OMJjDQE
trimEyzam8OGGlmjF78XU9JnDCf5fbWmOixgZzRLT0+S9meGmfGqOtBWEWkdoakriT399jaGhrRY
UybTRH3jFEHaiNRFW/tuwhmEASvKb7dVulIGGXUlXKsVJLujURCt752AIdf2dJX9lWnWFUSSIxUu
7qEAzCspX9Op4PcEbP5ir/jDVzXfO9rTTlXYoOAkPVaXAohiWIfJU2ujAmIGz1K+R3T3BZpxw0cW
HI83/zZEFTFZIT/tNpUmBRktp3LN1cz+73+q1ptIPwNm5zLTndssbtEUSpLpUnC3NryQrENDhtxr
omXr2wLgQFf9bc8chO/1jB1C0XgKBaQLcdmOfzfFhZOWVGmlUB006N2p6lRdjRDnWEYTx1oL1Ehy
75hnu7/hdtwBRRWAjUzoeO5m9QMI7yMogBECgzUYLQSlDFxQyx9nKFrGKo4NqfPJv9qJRuXvzwYi
Xp+YkAyJcq39AA1ilcQ7I8kIU7NKZ/Oe7Hfbm61vWs5E/THZ5Kmhf+Lro3Eakta4N3tdr2xLJBzt
XItgEDXyzHcVW6dg3Xb11VUXhfBXaxy2ZIzlY7ax8/HB+bZofzgp57WE0MRjKKUSMx/6xWlCZH01
YFPdYQbvdm2eZoWA3uLykcTI9/iaPX0tZ4r2uGkIkrL+GEFZ0gTnxXcW4sZlJL/ve07XGg3v8WKz
PtiEXgz6vNhu1FDi8jXe9R8yZvN+pdU+ETL38JJFwp4h2DCpc3vHElkhjDGEk7FJAogZXhK0wkly
zJUxr7FPWOTkTQ+BC8IYj6B70fjKCcSSHPNx7WVAU87xEEQGd0qnPmYKZCWLmmqN/vej3m2lUlEC
9laqFtfFcC8yT9X7aY40GA9tM9JStsP43hg/kLsLuGAfP83qx3Ib2FH2CdLXQmzWwY7HBT/N5GCc
aQPTR7S51zpOBr5ElWZCpHQB86V6pQpFp5xBUfwbspeq8cOkhmZCXZo/YBwewLyn4wxZf1Areo2S
ZHFO/tzx1BCjaigcQJD/12Mhl9qpZ8FHtRShUE0IOApndXePzV71xdrRzymCN7m8GmuLttjBkyAd
Ej1veHtnkddKrVNjnAN9VQWe0x9DcThfg4AfJiYtPibTyYHQcw/cMY/d8T8odPnOQ2DTyjwf9G9a
mpcju8pfiwK0hc7aGEy7D58NNkIdcVM4QDd9o1EC1C2tej+WFNosh/erumwH+gHls94hNhEE/6g/
IVpGMcvQtXabJiKPRxPebj4oqNXb/xHp7cKk/B9nAZ6Xd0TWC9lvbMleSERonCkvw507rhCvvE9h
HfNQjbdL1GhrZG2bn0RkI0YQCI+yuz7tHrxsAui8cZPEul3dLCNRfPBnxycAI7hJOLpF4NXq9IhA
W5i2rIl5uaSOu3tmtDqntJxtuPZDTcFW9lSUXISkYjNwzAC2LucZK76KXrS5OkyD7dN6we1FbDKL
z6dEwENGGfN8azYflv5aqSrCZ5mVZ3o7b1nueRHgX1937z43PpGcUAKKUY2UOqOVeXX7OqKFaBq6
n63aY+pEXPgaqTTt1wDX1Jd6X+undim9R7rGgWGlAMBCZ+8tSzlxP6PoOHFdu12hVNAfVqZeJlsw
qOZqKSF3aazFICzLW2sQgqoB962ScyMM9uBGrMOlZL1d7lh2ZjKit8ZDCE+85uzqsV8gxmyvQhxY
nwGNp5/HJ+ulAJYPGxbHdoG7UZDAdyoaxU4c6VCJdkscHr0OX+0aZT7Afg/hbSIkB1+XKWg7eIra
L2EvZ6eq4gPUdo6rEznCBWD3G/qQZ6c6qNU0WU9y0A+EvNsACBbrcMpatjLC2E3/l2Jjt1t68exC
y3835aOriopPCwSHtfZyCNU8vO3/vGAIwNxnK/Gbza6MJ3luHPCJq+Qii4dTW/vWy8QoU+b2Om4c
KT6TpnvzR9QAoQbTNIX/1NWPlPE9Cv5pSLGO8YTqZ33B9sfDE/Ttp64k+u0ExF7igGO9Hpcvcf8W
p6fkSHjAE3CaRVKWTble/h7BqPjoB7MpNHzGDEDCv7QJ/IaTP5v18w5KVdLL9PN9o8D7Otw2S/T9
tuwdYA9kx/bjJmeAyAeg79I4HSU9GNvUcHmSeDWQ38WIpJK3f7086bmVkiwGy9lpToOdokiu0xvn
objJ4mkl9q2XdtW2/UAZUGd3EFpRQM+m/w990FvQI3//bZn+WnoSeu2+FPu5/++VdyuuoZ7YN6Qx
k07oQrkzL11H2pt6uz7mR24i8evvCiLiD1XTYdiVt4sbVCaCWtavix+8HBiuzfTQOvUqYFOLz9jY
cD3hs2fhR2c5jkfh0d1/mk8EkkV31+Wu5G/PzZ6nNqhmFlm6HCLOfbX2M8v5onswUWVWS7rxEvN4
ArVW/CzVbl8M207P/dzviBO/U+o57BvQNbE+3NM36EqTVUPtEhdqn4TSMkf4QGUXJjp8tGhw5aBy
CaSRn8bp2WxUDY/k/53rzxgwiQYQem936FG8B0Jcc0laGzEldtAENzAHGEdcOpTkf6nQxXLV8wiR
WKu9EeWlCdU1UmgjnJg2Npwotr+97FvzUP/SnPcndkSHx4AMQiZwEIPu7ZopOE94LGOXtr+CnF/6
Dq5vIPTkWT51dIUHpG6ahOdqnGvoN0sf2tXGR9dJNEbpN8idg9QVfUiSgxgOHWpdOdggV+KfLaSn
wxg36asiaE5/pwIMO/D1Xg5B9MMF82RH9duEb/tSTcm/XpbtitHn53jbvgl8WoKdrG5b7E2VuV5P
yLA6J/bPATKflFsNdQZKfnGdQhbR9vn3DBc7SMZSwthVlDPMD6+WSgsoHqC99Sf+uvZ9uYSllvFi
Uz/NLpbc5ahUTz7tvXnFH05Z5Cw5mmKZz83sV++eHntY7/EsuLEUWhnezHnY+TGUfbUQs9UDI2qY
3XGRQUQYkY9SSYwhqEaXGpSk40MykAQaWM3p7lV0xwGj9pm8+wqPfik1NZy07ssOSis/v73BHzck
H50bjocNYLq09Nj5mpPpAwX7VvPu0PC4yQUsefg8ai/MP3zscWNeVNVZNGWJDtDW7xljwmIfHafA
NZEtE7B7eytEpVKry+pOoY1JtfJbt2+somBEhADoEgRFyKVOrVBaHIGsFTsErvpWgXIidcBv87V3
wNiWe6Eg1k8EqrmOcyOWFpa832cpP+M3JsACybnDPb8rPj54zn/lISJLxFCZaWc2CZS1oZQKqxNJ
Q9Gme8CaDKbLqez6HkFF9CXo5xukLqkBpm3wFxv2u1dw9CI/9CdD9zzpBGky33v/2h0QrXVmor34
sGhrgyIZkUeLqQrFGim60yF2EUkjxoXt/qGfzoFQY2GAjED0j6PtXMwApQYvqHyjKtgZSHrV0uu/
OwRuwDIVyT62+y6yXmFf0LkLnqKCRwZ0FOAHZHxLNei/z8JaVAfi3BTBZUVb0QQ3xQ533hBkSoDc
vwPgxprkjDXHJCu268UNHzbwHDXN9BNKO4ibYsIruAo1i97wEZf3dqJpoushwSsTjcU3ttsFVQaH
Lh5eZRjiA3m0FYakxtYpkxlIxnyjDuUX5prv4Jf9ASu+W/XngLd5mfUODWi1P72AiIs2LVuYKJlO
T+RfHcX8CZ4k2xW1OvJRbAlfamcpxQyTKLYLPZIBFNi1aJPqlSQuI984Y6GNGnB2X0x1cyrBxF7C
IFJr3Dp5We9zsYlMyxFV92IMLO3Z4EyL31+KZetpTsw64OgAkAx+G1+IuNtuNN4h+9LiZwflWmrg
X8PNt/BKk7inAw/yKmqUGzGtqdmX/cKQDZ7iAekJu8a3yW7zYgqdiPco/FIUk7B/lnF2z/XTTlnw
5CSW6rGgh6rFxGfT0GvZr1ysqTtp0sJV5AO1/h2j97q+3SW0QPVdBW9Ssh7TzpFTBOqEAKrmlTVu
oTjxJTxtsaJpdTltHhgS6LfXQW9OFiLHA/D72tlqPRKhe0kAEcmwLIYRIMJ2+tKFSlMlyp9fmPKl
zNrvUXcNxO4st9uT0bKiC5zDvE0f2FCW0j+jZDOyuKXwFipNdF9O+wi0U1jQtxg5jXqip80HpieY
JTpqHp9WNA3PU3bHHX8At4A858BEk3os5BbZ9aOKNMSgdSAthwFCG9ie/AuVWThFHbaoMHofM/NT
oLhcHjlN37FDvvsXiHLki+ofg6ZiVOQgtxdtwybpnvP+FpQP6ttVSOuMUzcZSOXrf0HMLSZv4JWY
u8v78cG8BQmpm1X7cg6IyAKCBi+hY8ip8hf3Hheh9E8W7zjJIKvMGGEAkvsZS7dY0G5Wshm0SAHS
u3CfBat8LiGfFWQ+dTDFXY2YZYqoROctkXIrw61UxUVSiMTfGJv0tcorn6la1eyszVoQqKbY6yI0
uufTbPx7+iAxzB019l6776M95AUtKtPG6C9whZoIt/Gr8gpYq/9a/vieeWPHPr6/c8fd5IK4Jhr2
d/OomKhsO1s4bwSVseYtjajKD7dLBMng1DIV+Hs395NYEKIUfQ1CEIPWAKiQbcQm7l+0MYyXrWlX
VUO5ixr5bGVmO+gYQlDOIXAcpJRE7JwpDiKYvsbJxZU+EQ4XBHzwm0qVxzc4AAeSc4zkgseTIWLA
AcESYYJ5Fizje2I5pgUOZFmkmW5voxGyDtoY03+kggUxrs9g1Fgh6yShc6y+MG9G4dpHllXxb94E
Fyb+OwL6KVwkS0fM24gOucM+KReb4crDihIjvfm0nTvpTOe5sumkg1SXjhWpRa1YKpye7VS0Ph4g
w/BRt3qJoH4djU598HYhmCAX+H67RaZ4/NxEbhOlNVFmzabzuNq4ISpo5/n/BsIaesyZXYgCvIVq
EF7RsRBUYPT3XlKbDQHEKDa/0x75/iipvbvn8Iz8VJShnDi86TrFOOUN+e7Ws5lm+VQ92Uer3g6o
6Ztj6BlSRDv47gIFu8D7t6Di6TCge4A0wwvvNwU+fumgjGgyDmWIfFbeofA37U+trx4TcpHYt6g8
tFaT1PgSkQDMDh9HWUc0x4VRCt3d9JDEXc1yBQEoVT72eQYnS2geIskcbZ5LpxNEVvPbbwPPZBN5
Osuhyc9k9osnMcNViifFYmNH+vX9TtO43q7wH0h5B7wN6XGCUqzauXc47Z+Aq+Ww+fyorYATiAEF
W3e2vkYG9B/SB3k1bqhdfMho1xMLCWMUikSTj2TlCfP9Ce9uHlSht+pF/fHue3HKz4jKzUtIIlNm
N+0/ewUd4dQxvYUWsCc7Fwbo3i7i+sSwnCw2qMdjWHp8BA9/eomS4BnUNoW7S/8uKzXmivNsCjcU
kkck47dmmEtj8rD8LQKmwZv0mqIixTgXHno/j6gwjk4tef1ddaiX+xloxXt8OgUmFg+0Z+7LRsmn
ef7bzPkEufCyxj+AI6Srt0LyH6PbOt085Ki9O+Km8QqhhVruTZFsu5yuGI0nBOemrgdoDzH9Nfy+
PPxICHIrKV1QwEgDoiqCBvL3pJccrDs30hJrpDUMcmBEeH1UwkFGbh+O0bTXyS78GFUvkh4JG8pk
Wd/t6QtmE7tlMJlF+ULCEpxj3+dJDrTu7/KnFj+QETtoAIj8Vaiw5+iY69C1UvpEQ67j/cpcZMj6
qalU++6+20k3dw9lHJaauGxTmeqgJ9r9EFYbMPya6XLqsswjbC8Fk1zHjUPVqJU7G7Dxhq9LKPDo
8xKMZf0EwGC7o81aqgx3A6mf+YXBXa2AdoUZVDfhFzZqL4rSRVIB7rotudPabLrDf6LauQR5x++h
+HZLlEeClNxy6m55/jDFycQ9NguVMcKxWo5pLQ0OHtB9xFgopP3WZXV3fX9CgghE/W2wWNY8jnol
O4t/OEAbmQrB2Adzijjq319oCL3z1/lH7/xhO0Fp9rRWkaJu0uK4Yjj2HfaOD7tNjNqH9uvSIGlf
TmUsvhNZNnDjw54MilES98EqC/+/eydoFxZvKdJbzWj1Zron7k9mslOhsadIAVRa9b7+pJRZiGva
Hspx0Bz6e1BzNjDoEEbLcljglqxu942FCMD3B4RwbusuLVN8/1xw3AHna7uQA1dLSAHagUvDrRCR
3u2em3XjohBQBrCmYtN7STKjFu1H5QfljA/BwUkI0L6gXHnJ97N0z0eGiMYT+0Kpi0XSHXKntbSu
BRMjHIKW2KX8me9Ekrt7DYn1GIw411IhPigAUHBBI88zeOcPkoaAfA7u5As7aUcsKlL4M0dVLjiq
cdZ3nnlQi0bOlLNDyh+pWAIbawy9m7pFmvXv03z3El2bdM5gXqY0fmrlJGWtJ2t85v34ROEhAywM
5nO/5awpN2oHT+4FwGEEz6QxE2bfpEQ9iJ5l9bXjc2hp2XpVxMjPkgBhRnthZAXFiaZ/6XwWRf5K
rhjTayM+dCG1t9TTWuheKCTem57kDAs80Msg2Ar8r9pC7KT6O6fblTsNIRM8q/o0PnvzbKEABkIh
nhtX/9lghk5Q2XUEYeHkfuoT463p753/i90Aj9Juabh9J/uWZQj/FZJ3OuVOo4GkAfCihAEO2GnZ
SPON0i3Wub1BlPw5att+CYzTD2ABI8TGmxxV06FvYFAJtjvHls81aRvDoUToyRF9EL/SbXMyWtlE
dzCNfUuY5LL0YoRK+mmIcDCCEK8438qlp51BYLrUk7qDafw+fw9+PVuLrEANST+Oh8ZOtOKZ40an
Agvu13ODj2ODScAMWCbO3QZVIVoQn8x9PM+mN/f1g03xiYT0jKXGyandRVDJqScmf5wUQR4zYv6F
NK0eY0RouEU1Dh1EoxwKwhKx9K1UKkuJojsxZ1xb3kNCb3TB3B3WcsqsgPm5qEhsx2NcWh0BuZV+
Fx3BhCeIfuX2MVjnQrBRCqxWILoo0ZQM52H40wUj6QT/qmMGNIbbhXOR/m7R446kJT9aFepZmfp0
/YrLJrHU2eXLqyp+PmH9lLDegZrOy8RiM/wzg6EFOM2VZDgDb7MH40OJy9Epz0r3VbxGbI6BWjtQ
EA2OTUdcT7iTxOsVAj8QIfj5nZ+zi88aI0U0QO2IO0eBycIDEQS+lSBrK7Gu1t2B6TTeygZRjgKJ
PgIAUjJRt4y90XvYF0LQvFuJOMUTmCZY6eWGa5fwM/oIyzgWvDAkyqc6H+moW7SMy6GNfna6Xc2V
ueoqxRwZX40LvJT5BTJBgvnq9QZW7nIwQmDiHCypT0G6q1c5zSt/DtIaSsNTKStD6COlRJ0KxB/B
xBf3dDAIOSEsNM2RnITu69WxnEqc+kFgMzl627ZT0TaF+kQ4Q56omW4RwvhjirbnJHqZpN/ENLyI
1YjlAiY/ufDld+eFUPbQ2gSNv6NZ4YPebFSC/LWC2KTEpnB48eRHLKeBtCog2NYJs/e6MPkyCiXd
NSAwxGDnsmoP88OsqC4nwHYPYmxNJVNlssOXM5vRw9eFRpvJw1ES9RrQXYKpdyL3I/nmC935j2Y/
pAnPHgO5KgAhuFmgBxuKEHt40IINwZsdEc66zYFA3Sz2WWzFOrwhYm+MDWM9DTXpSpg2YbBXGHau
v8tlnc8SGnmMmtcH5OXjZ+/AUmTKxTcv1Wapf02Ak6pHSj9SuUrxPTmGoDLWbsGOW1AqE31P5P+y
cM/gYbDvwRwvm/hJhzmb2+uZUdmXe8ePArk5j8Fb0/sBopUxvABEsZ+1Zg3fAxCV+FSSFe0hEGtF
ulsc4JIJ6znaqSJU072nsqJRPKafwdHWjtwehIArunKU7dv2+EvGsCb+MK2PoOmEXvi1pl7xLk6e
wJGxfdD9x3ATQkxRxbCBtm/kKHSVZ14E26Y1IIuzP6MNiip5jdo2vCFFwXmkHVE9WvEcVn2x2tdV
l1zAUST0jk2O9SI+KY24vJ+qnRVF8L64VAa9Klc3fByHhFLI1Z1ETvbN9JSzwKjjYc1caTy/C+Uc
p0mGxRXrGVfJXNWTzAhfMzrq184V/EgWRxO3PHM9xo8K85sORWltPNwsb7EiNpA5kFKCuGD1z9jQ
4Ep1bpTmK7odGUFgdLQXVKGA0RDewzrO1c70uTnSjaJMHmrLSQAvXtX+7MZJuW81OC5Iqh/pAL/b
AZbLc8cevzvkyEPWeWJM3RYpwM5Hg49KLrF3dJRaBIbA9m69xZwJn6UcNWreBZqJQtmVPhXwv/4Y
BKD5f8m1mG71Fv6gl7nz6iWTmRCd23s2O/V203FTs27Wk/iAk0hQ0jCiT50pvGr02xG7Sk0VD+RQ
rzHqBiUwRIUsV3u1bK5ceJmXKNF302loruI8Z4ZruDQq+KG41gse2GvtWLKG/uuwfXBvpSmp6ylo
XagsCZ9GvZBkmIG95jNs7GYdLBBdCIPc45jM4ZoTwKDtmFxHSZ/MBE6Rvc4HFY7f+GISMGNIU7T2
8GNu3Stqz79jEbReXELwq221g5comRD6QuqON2w1ObJIeghluqtJVdmr/cop8Zqpe9wG1Pq1kWyl
fd7UasHyCce+hRW9SCsjH17zxV0SWCr68jATTIv8ExttlTYRZbOLSbFvg/l+u8tNv1liTTjl5MvH
Hv40pRNC3IywWHiRpStb+mcZAbflUH70F05BZo5JIPhyP4NZfeMll0zpnMYOjRaxZ9wKquVIyCVp
EslJv50izKdWZwMx/TXjb/CSDBEveAPDkndU5f9h2paBUBBhlFTrVLo2T23pXlQCb2OIe4J6MWju
n2AcA/QdXLWW9bJwY+UDQRp623xiBpXYTJV+3+v/hnrCvJngqpv9/In1XdwobT+mIP6/ySinhFL7
i2W/h4ALkTKO1BhjmOLF6wJRzDIRBcxuhUfPjuWb793J1kkaE/R4OnfrH53dxjUCqGvng5sa6RxO
B32ML0HE4fWmYXywXZQHkyMNaZTLMpJamnd95GiLintOhMlqh/R2uBHOs/ZjgrfimHLFwPimLFRW
CTFEHyNL3oQdegc7HSMssdEXIFke+qJMxJf7yMjnNa5fZv4uoSd5zS+xADWEBjP0aWWahthj8m4W
tKnR9N2GLcJMwrcsow7RYz46IhUH9XHUxUv+iICqUlZIMTiz/asnk3sV6XtC8APXmPUO7o/YvSnG
xUrb9HGj6K4mDHxm0R9dVH91MmV3XyO5dseIWoob/5KZS4JMeTpm6JainzyO7C5B+BFJTiFAUgki
sr1c+9ofUSnaps/NjS1cpez80357WbiFl31bHaxqYcU3f5E7hJJqgijSWf2PBYWBAfzbxPgwQFdZ
7+y90OQ3e1qv0wiVwTQ+TCJND/NOug9THTepg1sXfHfzgfQiIG19hwj18XsBYfI1Ug2QzSiuuf/P
NWMZWts8zcJd39cNHCrGmoEt7StXeAaSM74gfdJWccOdCQ8IAWrvXNfcdhy5KuxYd2KV6FuFoBJD
bBF/bgGg89KzNUepRS9OxMXeEw5qfZRSWrzKXm8Cjc047uxpha0127X3JMtmD6kjpfbZEVZydHnN
HK1shTPB/PhEjHdZGeirgp+7FA0t0mk/vDeQOY8PREkPuBsU/v3Qlod5kmSjD9Px39Fxo6ttIEbx
S8NSgTk0VzL+rCsYSVlOrimFKMKKmPCnzUfJOHtsA2XnNrJCAqdoLt6CBsb50LMw+0hWcf5ECFzE
7Fu7LDrpoO4p/gVH03sZiQn0AFLtTN+M7cNomACFEJ3U3AcvbEWOcevjnJ43qQ4fqAV3yUkK5jm5
C22xI46+rbZW9vsbt8goqnuavdhI49yxtco+NMz3iODciM3e+MpBkkeBJQbtRYAbVI+nuMyV7lQs
7HIxf0qlsaleIT7iH7YNXihiSbBkNUFV2WaQUmxGU1dfHl8YEQUly0y/aZrs0xhIJ4YeA4JKPYqh
Ad/ZzlbLHE0WgFddp8rds07+V98WbcqPhOUYj9cPu8bKIVRHgpk8YIIe6KeqxAhisCVqjET0v1qt
A3z5dFw+vtlvmfJrZYMP6UsmKKas91bULjtlbfJ8NHkFWda/a1maoQxf2//9av3YMyhRVshqoH1e
alV2u2Ylmn1OPeqkztd2cTAYOzGxHkyK9ZBZ9ysqzvaHVMm7QIz2N/OAUWPUtSLybgIOecMmdeuC
+noV4M3cJZlhRFpDkV85nEJ3aDF/a6tNBGyuUg8zDTCrP3JvYVpNcxqroems2grTMrcklxZz96Dv
WndD2f+SUUNQ+1ElMQN0qX41TVUm3dA9GgIqYsjaLxDeLoiRSgbXNgqomLpM6tjYpY8CTQRadPrz
USLlouWtcibLvsn7GhlYxR36UDNome4SBabRrwj9of6S1BSePwaFdKKirQ0PhHaljrmQydh8STHc
rWtDcS4bJe4ynszxPOqBDxDoBBPhHNx9IjOkSvJn+yvQlOnHSmMXqbRYOO2/OxfcXM07QMPSLof2
mpcZ9Bo4ZYDmvq/5sG2GYCOtItkEGIAU3kS4iXv83DVSdVoKp7mY/58O90/tO3HY3D0OP9V218sv
6l5vnO5WhLi9N/lgB93dZpPiA+43SHIEXLRx27BRaZHnEP2SsoNI7DcM4y/WpkjF+6jDYl5HiE/+
p7oKXPNzab2wbePk+Umfo4Lb+ngnjcW0j3OhinwKW3aDY0eQmAt6/Wbv8s+N3StXhdx+FfWGUq3O
k2G86j1ftpRJNjMlEb5WlnILNQ0ax2Xkd2JQNgcbfFFXzzpJU8ep3AEcntFYBQiiSr/wXN6C5+Mp
/XTuUQqUx5g8GmQtLq6U4aEA4m62hF7TzXe7oClsZTarWsGSHklqlfj3GyAW4xYdINOJl8X/CLnU
/epNXVp0mWRKFCJmrrgMvXeZW5lVxiRTc+KqpH6Uar8Q7FaaZ8VoHOZ2xYiZsyES4X2PcpQANRBL
F8y2Kpvhw8CQ6ao3YUhExfAvbWTOwajoRaY3LMIvLv5QGmBuD1MdO9AjYpBDaIOzBdikAShjlrmZ
c/oYcv0l19YeO//nhSs6HhVmYSTIvTqambZtJPLrKTbGfOvd/doTk2w9LH57eu0tepPAV922XOHd
sf1lzoBqbgxTPpVyvBWy24IZiIuv2rSGojlvZKc7iUaBnYDdqouRm+m7UT4hhn1lSMb3u9rpCej+
DU8QCHc3kiEMGuFrCcSTMBOVZiO3zgb6x/51LqNrcE0xLpaRnLkiv9uSPSTOw7Lv60FKawYeTjX0
mR1zRZA0QhlutRe5HHIzL2YhHdQ9jLF3iYvVsK1Sd30AneBPAhA2eEBrcK2JMFWMhEZAaQroxKao
H8n/webSQY0nOL7L9m5/1ns3/Zn5Q1pFHKW3Bk8lzAVMKIpVNN+wzpSZKjV663K5l/IUkja+To73
njGJmDj8SHB3jUTPBR7F7A51NGCww3yXErm9UH9g//EC0Gbw0g+UhHTTwQSvg7Jpk9lfAWKHevQ8
UDRvRmsA+m/5wKClDjCtRDhBbI8ltX0cei3xFQLJQ2jqcezmI1t88KSfj4ICA4/+JGtkbdOLGYpR
zg0b6Ubw3ct3PVrQLRTbL/69Pz3qLu6plKtcLFA7QOcwidOtGHbho7+bztfmGXux4c80VvImqnDe
t+P3tQ8WmTuCIkK/tM7E+QfeWtUF8dDSbIg9wBcwQUR21bk8zRtMBlKesgNO4uFeKOOpbxGIUQml
VXmwS10STgcZKEXIGbuJfoKCxNZcfDf2ywoIvwShcKEgt95Xk28/ZvK66ZXoBPkbbBCpeEcs60wD
0qr4MbmY6jq4MwRgNw5GTpHG4Qk9gsUzzGfY7Lq+G5MwO61Il6TmJAyOJ4d40b4p3Tsuvy0tu46k
9mqLEZl8BBLP8YMdibbvhfS+LCrLh+8gyGV0O3YXStjZOs9VgCVHHHFywdXAup8VcIxIl+teVspB
sxtbVQfP2UfIyMJ2OwPI0Cx7qsYygZPAj2etRrabgMZnpGAnjXautD4moTXNYiAuPoZotSAPEchh
rPA+9pGfdd8MpPTxs4iAKXSnC8BbmKXkZoXxzxVzLnU/7U+L9krwWPr+ZbxIbGz0/X3SiFPjz9Z+
0fIt0HVQ80gAeT4A/WwgVQlAxT9TrKYm+EJskO/jEAfJLIg7FQQnYalSHtQCi7AVSDoDEUs7A65M
PH30v5Q6d9LRC8WKcr91/w0b1QHopphrTHtrTaMPn3uabbe2/Zb5wES/fmIDuOzgDaVO1nDHcCDk
eW6l4IxkLVn34EMJaRUdFcrlGDDrUz4kHMtY3Z1hmg3Gq0rFGOf4u50TWkwfZuyRqk0QgSQjUy0c
eASo6JozqYK0HlBUjqbbI/ykfFM4bSso8skzTmCqM5b5s68N6DQCiL8R8+RYEDChz4AMCKM99NZq
eZyllNVuJydNltFqKLlqI2xVUouP2Y3T+sSS5jsW31m3SN1YdpUqSxznfIbESMmEuD+agmy8maDi
MDgOoP1BCt866fYT7XqIfChP2aj1smOQxLuN9JtGKSE1z79irvjiTVmCGc1noalkEfyfqJSpRlqj
a2yxmbyiVSIdMvV4NNuN9Vx/ET+au1RpCbiSarWkHLoeCjxXSYhfXqdmiclVWZa9aJ332UNl+XGf
bVJEEM2teo+txMBfRRJZCSUR5+pskXwPb8vuIrO8iuqdsiIAPR3bJykYhfm9RK+Ew7KlsrUYlxOf
ehnW2zXlM9EH10M+Nq9rp9a8YJLcNz+1U6l/Gvd00FVvBwLI0QXG/rfVqrQj6ANcP/wgXhZYb9Wz
yeiv8uwaaQdl6aV/2qJ6xXQ7yH7NgA/eer1FlZItmhhHagt3JFHcPelq7rYPHcxytfD/MQ1LBX3F
MgD0AjRo3UQQsQrnF0wvcpfy+9xeWvwEINIbfG5xXdF2EMvPsfSUUmBQ7B+GyqqH/4GBdEB/eiKG
IAvuxFRpjwoZkqBEK6VTNDfkGFtYHXuWRQz3QnakB6bzaffQC4WV45uXUKQlvG4EHQ9eH0ylOVpc
fftcvq3ZkxoLlz8T4EUm+3fGRzEee82FZs47RvWCC6SfiSeAjt7o+rYWdQ+E2Zq57qEsEOdAs8QD
P1UWT+4iC2JO0r6ZBe4cjwA4fu6PRZ/mP50bU8uhmMv7FmRJjf6vDKKs5QJYWWp888j3AkOppzIL
o1UgAHT/CyiZSLPU3nKW4WLcYa/HZW1slZZpDzKj0ytaxXnrZz8uOBJyvXRjacgAs/8wdraP/zZ9
pAC9h3mFLw+X4THiVvWcbCbGUjvSuLlGzFEjebrC30VoKTv3g+2UsGG8DdYna+7ent7EaOGeJtEl
BqA53EvcXTU7MNSBFrXfUvQEOHBK4QdWSCpIOt/uyDv4onAcey9ycu1haxHj+1fzz2YQD8ta96b9
YQifRE9c+uRNWKLdl09W9b2wCe5b3mVQHB9xo8EyPV84s+bOv2hvt+pljQEzt2038nfw8stvQ0xi
y7qb+8uTN+ah2ePf3/iyreMUBnrk/AxcdxBeS2NzkZdEV7cVBTd4hBbCSZZG7W/z64b7fpCIT/Hg
3Kl1qKUuCsiMU4UGZPuo07BajNiEHjrDpIZTnbzzk8xzhnXtKQ6uI5+T1BP3NSSO7vBJwn298WhP
J27ujgT6DLxwGne5UQ60xYNhA2HSalrVESDd0o6p8KmRKEK4tQM7jh5wfkFg7bV3avjX7zSpaBjF
2bpJXmox0Lmwrn8wUF6M5cyULP+vXBXmaHqfUoGCKmMRzPTryg5IQeAwZvxmdSqIyJXaEPLi6qpm
9ev7w6bvBc7Mlgrz+N/fo1MBmTWxHhj6MOYjKjnPq0/2EOlr2sg+VH5432AvSCaRXPWGUCxIASju
DRabc6vqU/ofec19ceZZHjLBWqzM+2ZNyRiNh023aBOG8jexoM8/IqQaPiCAl0WM8sCto7/c89qy
1k2yatybn1UD3ioy0qYMZYfXGV6euJm2pqQEnAN/B20gI3VFHHpnW3k4g01lMiQTC3so1OcHi6ZP
WyqeyLErNxLK2toe2AkfjapjUmSf7OACSnXjVVp2FfZyd90g6yg7DtScGBi5Yv3Mr/82ZiTiJ3wQ
t6ixN9PQkZQ5MhPz44NAanADjNaXpTvUVzRzxYL9ftw/nVQblUWkWzuUHxkJQzN4BBHUBsNMmCXi
7yF4d9IZi0phrptI+xDutb8AjqtSiUAHYqo/pdrc2bAw8ZNpJKzGMJOu8K8AKUswmmPI8O/rxsQD
oBmsYfggLDqLkhtejUIeyzvrMPF4JXc6bPAuAeIenJgutEDP5SONsoWxkFutFmS4V9OhHi3O8eOK
oBDaKCTBhz/LXvmz4c7n9du5aTHca/mJaqJ+lRg9MiCgUJhPVejY8I33n2olg+c0hOOFwqC/ZVha
hCndT/dzX1TL83qktaUe+/E0MTEZdGkzQE2ohUC8P6SAHTYy70k8aV6m5u9RqocllNF0Uj3keIZg
W8IxNI/GxNHyLzGAYtUrxZDgzUHyVhDO0ceZJDYEfENaYqr7qOTM6CaRMGeub+gq+pvBmMvqCSGv
44oWJCUjzMuVWV0RoJtSGlO3/PSCoJDq1Ppni51p194VUGluEgHw1Whj6btNBRP40eULdntITXTn
+wxvpygK5udK4tchinPTGU2VRUpcQ8koOoRUemYPBo4SFTHirYZbBY3QJiEXJi7qoe57T5Xbpv5c
QQ+3+4YkBzAtTg8d4IJ4BVWDfv8VgMhS43S9O/vEkOGqW+B3zTD+NUfqVjOZuZUQTPwv4MB2Frnw
GlKD1LRnOEncEVQkk3BCg51Bdi+zL9vUk9JqD+rOBiR6odGjoZZI0CvketziItCDumXXXZP5EDJ4
kWW+9Egk54/itywZEZhYxo8zAMz+kYpcs7JP8UEWQ8o8j+pKFUesR2GH6mw15gatAQ6TCJ+3Mnk+
lP0Wgmvl5ftCKSrNNx22Ve6U8M5lIelJsMuIM5S4B8Y8RKHIxTWEiISs4VlnCbScqpfZ6xtVRun0
MadsdDiBRn4uS0OLhmuo2PHRuswH1TT6N0fHakT3spAGxD4/syYm3mj6+N2BqYBBCYfzYcz8XuA/
9D/9Bnn7qYUDJhbuywxykrzoepxUt8ShU0ihi0fKuFf7bgyva7CMC0qraZ3tnoYWLuNkr/aq1WiT
sLiZAjJyyoZ1HfTvF39nUmQk9oL9qiTuy9amjRy5QXdS7B9RakL7LwRln8ZkbDzycCNrCbGZAWrI
7SRL2jgMiazD2X0/JaxUcR7IXyj+lN9avsAbwVCqgO4R+WZxV0sAgYGZWcTTjtjLvvlyUn8iBC+t
LA/rKcxJAafq/251dxEOtEeT3Y79poDhe3LohKoLfB1irjeNPx/4grb4XMkPKWJZAso064xfcHdY
+PhUMwsti2PyT2iFtXVLAqB9GzNiLfYD58fQtdtucAr55wKpfA7fo78mscHs8xM4w2Oh8AGh+Cte
9t7GUXnyBUVcEkyEkhS0nrCirPV2nnz78ZLbnDJHS4Ylw17JGcKHvS4E0hwpa+v+b2XtV8raQwb+
jqcrvQ7FmFfxSlUYFSrQWqgaARuyxeCed1pGyaR3QSoQUY8jCyH8HnkkuZouQTpzfAkAzWmz8hUG
Pzh/WkKgLAmAcZtCgblxqJKnCJqD6sABnbKMouO9aOkEqJqQ4SErIEZF8YVYTTrUYfUc7fcMtJV3
jzWJIeCJdIFzrqxFZOoynBEank+8auymHjlTXZDMFW/MzKzyBSjCKu+CiER3KxDDbL/Hk/El4gG6
ses4aYNQVZaUAh2HCbLdw+3Pkun7ZAqHWNjckkVMM/LP/wtA4Dw1yZr/NeTqyiyooCMNoKs/kpa/
YPSRuFH0SPzLia92HQ+jHFJ4gOxVeL7Q9ySPoMEsDxqxzd6ed6vZuWBugON+y7v5U05oC2VXTlJv
QhfLav8tUmxh2jeTinvxYf9SVaz94IrvlOkUQdW2JOOaRTQufPUfKW2wcPdiOQzrSbl5FicValN0
kM04I3d2RZlgfTctSORIc3JQ0qeXSv8WUKccVcDL0xbm8xKHYgHy/qLmGt7jfaJ9WnWs7GBa73ky
edLG0EeSOo1vK7rNpagdpv6j1Q/JQ82RTtgiiPe6KONOaOJ7bEERxQZPJq4nJiKKgzhPJcoqWi8X
SPbvMJu0afz/bQ98o6h/eziymQyJsYRdnvw6KfQuUEiBt9aOO2WjYxkEi8oA0Lq8DAnRo+gMhAqE
PHbW0iDdp6uC95aeatzUrkUYooSmgsMiwFK30l9ZqoX0c6rskY/AP/dhaLRETFWyIXvzqTZ+olz4
QU0hWfHaSlT+tsp5N4q19UUO7J1I7XU3OoWaSDQc3A0X9Eo8derG8aNvNyrSWWSykgbjQ/HXnWIc
TS665PdRVsOwMQSv4Z2m8CfZ2qNeG8mTyE1obu7T/kJU2LMD5GndAobp67OzQUwp4KvGhpnDzVPy
2BU/tLHiZ4YODIoU9VurpkdDE4fxWcIMaCHnxDdK0PI2sjPhyUl4CTlVWoRiOoxg0BK3Xk/WHoh4
JIOJwlvPMZwG3ZeQ4FvnXRL/gJBhaft2zd3B4oq5aomEbuNq/4EtuZfjKl14+oaGInYdqLWWEc1p
nD8YVnW0Gqi6Z/uG8l4RPVuDyqdPXpGRLLx1TcQgMHHh2Fws+qs8gXlPOBUILt2vHGAIGOdCtD0J
Nq8m8zHHSviieFFZYwZV3/j6YBXcgkcfL3TJwyVr7KWEI6+/utbiTqkAnVBGoFabW5mSHVjMhkHx
ym1jKbeI06cFmdNPvOAg+6by7BR99wxu2H9PrSceSkT5fou0UG67UC9D8IzdI09xqrCB9I5ocU2+
NvljD1hKeL+DU+tXLgge8nwhsG516jg0sTDoK9qg7qK/SlL/9oUYTqhZKcD7qqZaDzQyIV2vV6Kd
ONVybetGNfOoDelQ7qdzA56rawqiJZR140Ukt6G57QNoKE52vRGJbSCAkJHIHSFFvTJP5Oq2D1Dw
5/YMPXRT4E080cWXVxJFGhLOtJ6XW0awMm5UE9KmVvYT8PGcvHGbxf2883qtBS4S843tTilRkBXX
3/zvEBYeEMwiFJp6ooZDmrrg9zbfF8X5TnCTagtpDOTaUXr0ouNIxjoAmzUsvyTdArBa1aOHNAtZ
wCxl+vVrbniIJ9JWN2bCg5J+7ijbGHdJo1Kxlkfu5/jmfpP+GamoaNEjhg10399ymfwizglzI4c/
8ayqjmhl9Kl0ZPHf+8IXte19uBcOGgnR/bPS7cGymNuNkZu/Zadu103x0T52kp/rjc6vwZzD+1rO
jFt5LBaRNm5Y6sK++ddLYJxDqOG4Eca1yoELFg+3RdV5KFe8hQ0Yh8XZEu6D3seaEzk0Xt8QysIf
Suw6ZO4UdoIIgkKdlkHH+bHQvGl85dYDwQ+jJwDTCHdanZWfo4AQ3bZTj58nF2HJBeOdxyuPxxXh
F7o6q+JEqmQ/9QU6lB4LRFgyA3VfWdkkZdgtI+nEWQDXg7A6y27tZk8ThMsl/VrxZX32HCsjoA5W
KGGVfglX0Ro3Zgt1QYvRfQ3qB8Yoa4mVUa8yGnTIA+B0eF7/+44beCfeO6eFz31iLp/dQOzbIOgT
yjyhgObSq8Wnehfb3+pjB0jXm8gabcp97afEUZ4P6J7JHkcusv8g7JWbv/zUweYtnzUeUrSeJkml
Do/zolrCUtkSAfVeLOAf421Lwzi14aSMvDzclBD4YXqejC8oAVWV89fJ24Cp3HIr4+kr+U+7IpsJ
KqNZwJDIa8wt4vaKLPI42a+ZRE0Ilf5Kav59iwmSEgMZQBMVvMi6XPz9h58RRHcVFDjOSdtgGn6G
lN/gh+ODaFsPWc7StWzeWybC2bfyxRZdrNTY71PYQ3bGNeU/kRlLqaZ7ovA1Y4Y8Ta4Y1fjYkrDX
GGqgDCKieUU3osoqml+1hR4odyqKb2+fXH0ur2fQhLtzFAV4Rvsq+0pLaLS1LTKeNEHakWpvZNzS
DtANTr74wbbhb2HALWEkYY0LnpwtTHv4Gq3kf/gcB+Vhm/d7Tg3GyJgczJnmnpqNalAf1jI7ZNdL
liD7WQBEzzrB6n8vfwQvVRgWpBHtI6Pb9n1b4RyyQSXlaz2NSEmYBN7FlvU2ZCwkRratvQ4XxyMv
kA/B7aUivH3BHXJnqFzsJ5B0ebV53zAW1/nTNGoJa0C+Pw/VL2619zuK9stIk1tjKO4gsqpC8sL1
9AJzWyeZS14HBCul9SDqU2AXvxXlZ5jxfhZimTL3XBZCm4yxBumzg3BhTGLk7ZIf6I2h9Eaza/MR
fv2kDToXivxejthJpp+S36AEQpfebPTF4Xdr81D+waMh1cKwHjoKvzYVl326eS7035MyjeknUguZ
VD/gs8doKM1GdP212+9/AsMXk6m2ap4aWCIkmxSeLL7Rr9zAumiHwFe4kXjetRQtiL1miwCIk88W
1qNuY8herLloBx8cTjL9yEtKee1wpsI09LP2X6XDphr2kTYx/CVXm4f4jDDtcAmxGZhrIO1dbvdm
7CNTnsi5i9UX3c6W9b5u1t09TXn8z20pzWtR0y2T22iJCTucSO7nPE3BG/5VXy9IEYkl5EmzeFK9
fCQaHWhA/vTNGHZ5POcuUX30lwiGPTkeXsU1bSidEqeQJQsv32Fn2usBI+LxBcxNZg726XRigEr7
uxy0ypEvgqafhMDVYXFETbYgIVrYQmA9UdDQt4BihxwtWYymMsxFzxFVn2gC5dZ5gRuJ5/zMt/ea
akvIFt1EzRihkwMp3xKn15YAXW0BPjbf1ETY/FWO2aRyN7UZ7e842RrkA1yoKoyLfAduZLtJ8Ynv
y5cIunuR2K+mMlhV5VxczcYYc04AHaTnv6gEuEZvD8MdMHFYemH/8GYVljWcBjVsY/V6pdvYFMxP
AI4V5cyu180osLpOFlG1Qh7ciZPHV7rkn+4aaPOiOH1SS57lpr+x88IOjFhCjnBmyR5Be8Hb6QE6
e47Sks+PZBq0+7t7UHoyb9bNDFavGCpPSpE3J65V+JoKSKya3gWcZnwD1qhOQDfw5aq7WqUVISnB
sqvYVzbPflPTHuaCpqyubhE4HoZaU4XX7PjBFofNzyIroylCqMGmpa/MhCIo9yhsaW08AIqI6Ujh
rflK5pS2QEOKzLJ1dyHAgVaabXbxJ0/DCksJGpktiKIaFoxJ/cnq2rtsOMEyB0cNJqiU0fL9Lxs2
FJVCW2ELGXEISRbzZjSEInyGavWZf4XlCcWTW9rRg+BL7Rs2+ka+c2QNFHaRuqYFxzu81QUnP4nE
63iRhvwfEAZk+x8mLYzxnjfcdjnIpfaAH9PLiK/+732ptAPko994A/KRuxrANhtfYVcJpbRDcKb9
rG0hU8pjt8Sg/VvFYUEzOhO0KyVGf/StTourAac6rIs0vX6sjpDdPwRPEUJ9AvmBtr9rE3qsEALZ
Hr8eTsyrK+2XIRW+iZHxR7Z0karLMabmVNwtaSfOz/Z+r83BeqUoXqAPDG+6/IXzJ6jSi8G216bT
gJJyWw/PWzmDOFP4Ga1XgqXvWtymAu+5tOzr1AXCBttzN4VCurF8QyECmBio/l+t3Z36EUkXjS5e
XtQk1xSA1ILfsxMryA1saCWgDuuXdbl0+y0UOGrJvdpHcp2Nre2oosslaSvXnGkYD2KmXeIbsVkR
Rm5tj7MpVOWLuWWeZyE3+kn0oDz4g+CmU+YE5o6vn0ShktUIJFRvkGUkW5KHnqz+e/zDNtN0Q3O9
Hf0mDQhvqS1IcRE37iMKokgABV1Qaqig6AYE/Ksy9Cc6DBtKWLcx15GfEu2iDmIagnRz5YNr3RkQ
jWj4rvCpcz5j6H1Qun2/Ivq6QC967Ap3tOLwullsmsk5Tdoj3MDktXwUQty2U9/vGHlrmSjCblyq
ClRojFX77zvmCvvQ7Z9Lg6cG3DUxs9oTQWYoOzNBJ+FVgLe4vhzB2FdQzFOCTjOlXf3xSM/Mtefc
lqkeSo1gAYRAmc2zrRqOKW+cKsp9gnz9L0TChSKRIw+zlwMogf/nzPUsaos19QNObHSQxuF/iBts
MCRVfKOVn34Hf3KMEz2ct4flxrn6za5Yfj4KBa0YtHAyfrMK6bZ/lgwtIyIO0zmWLf3xeioxGm8y
5kScZvNVqKUtPNPa5go6lmkccVNhZ+DQJFiIvdAmqAjlR1nET0YvxO2ioUp9bhcM/VhtsKdHKfR4
9Dr63s1w3jeKtg3iTXAsJPFhRh8hzyQoMqCG+UWUbXmODVxIjSJjMYSl2L3cv7hKmzm7EL6NOK42
+jWOISdtxj1/R7IA6cDFs+uem6oujgwFCGyAthTMKu7cGSiGWZTyETUm9UeS8576uvH/1u3K3bgV
7qHWVUB0g3ceb5PBUTpBV4xt7G8IUQ4Skw0JvnRNEk4p8TLzUSQ0xnxjkN5+L8lOsQJc6KXB/3pc
kagfXP6yZivQ100KitpVrh440RC8k5H8dPogUP9boPeBO3FlXBysz23gIIOgP5aMdOeS7ebysYiM
6gW0zUgHnxEXZqUJveU/+fpZTidPvKQMb2+zo5vMh9O1QTbzWU24bzf1fyImYwRGs7RIAUJZ5198
hHbFjAETYoYduhr2D1ecp307pvyAx4zoLYTJbmrZJC3d5ZdjKeRcKclV19Z2DRRiKftuQe/+gd7t
JFAlh3LnukBfPYZmsN1GIL1AsuXrUCU9XNVH9rzs47w5MXMTVaLHDvb1ciiHjS3lIXpBTQkut+jQ
EZ21cnKn9RPyNKHyRMzxX4t/yL7QwIpLtrZAu0NZf3m6S+rkMDlvuYBUssSEUv4pl0xkX8XoGeRw
LXny9yQGWa3Mv3lbnvUgE8PPdBFzpRl9yeJbK846QH18HfubalX9RNm9oC2OLpPL1QRnLe8QVygu
DbSkewan2Ue0LqyVFeJUdYeexfZ+RecGX/E/amv+7tSZvg0mTwXEDXRSUwDzH8TfvuRWK+TAHraj
eStztrzgZ9UKchlnAF353EoyLX9hHQXvsEKFVkd1LIYOej47k5WiXdoLeOzJ5F+FjLteubh3vHtX
FFYSRwGNggkP1CXvgq+vInuq54MDPEG0628Ktm8g0RWolNjQELHgDauPm8ED0mEN3bCAQgRVjVOP
ZLu6IZBVuaeNAygadR/132YN0Bkq9dar1wVqC4ajv60r++jSi0JejUIKtRcADHez8AtPSVCOfi5Y
fg3SbQAsbGu8O9/goFVpcTBXn29pK6hIZMGjoKhFxXO2BVb/a69I/hUBWyJnt8ZuR9BChmGC3yYV
YmsCJciYQfGDDPFzPmx8B9mWJCn8KDtLUYMNf9jeqTJ0gca6tPefMMURE+nQAOBoIBMjMn+VP3I6
TbYGUvQkedbXo9baJSn9NcqSRrSgW6CCAG5wNAVEcb8fPV3NxYw6cAG5g+h32Odmqpiyh0hIfp7r
W0yVtHT90MQgz8xHWupNjTWreBC47bly+kMxcKYP7+DSEN9LgSmGUxY+JfW1TS0G7DC4iwV7Bh5W
zxDQ1SlclxJI2DMWIOys7d3KYEGfGImsn0bNRI4kJIRDiGGcQD8g2lVMF9I/yRAv9P9qFrPshjVP
n9Wh+WUxaERaP5VCebkiFLGIPE0uVlyno/4wFTpRvfGeGakvblnSxG7jSfFRyOX4G7m2oGgJ40s+
FOZPUNdpbRCP+GXqpqXLK92tHCHP0rVvM8jYKphIWSne7rTn0psvDHL/qMdQ7S1Prk/jzi0NpIdc
T8iaRhhq1Rg9ZNt7be1Dh3O9auT88pggY0obw9BRQ4rHpe0NmlNke7fdoXutHH93OFFFSN8x8HP3
Gkfzhz4glKZ7dBxbqQIWUTlFbV7jod6o8T/LKZo8D4uWFcsEMyHNQmJUIvZBJZc7Fsx3POZQ+1lP
8zEEh55Yi273LhNjAtb1LGbLebQhriWzphfL6UUQUsoGnh92NMShMHVCytofuwIIIz8seVy4lV4G
woEFv7WolNRfXlsAmhpqv9oJRmDxK9d4YxU6XkJp/KtVSF4YgTn5F9bMnjDg41Eh9JpQghNtDvBY
c67Qs0A/IPCkBJXFVYvABBpVPJqLiC9+KD+YDnvSD8NDOIVSdsBXWjuVNbk0NIG8tD0HxbP7QIBz
zkL2W6oD2zssKvlEU2Q7pzmLkkZRIY98XbGFuF5ZZyosOFSZixDa0Vte5KJ+SUeAjoPLPRm8meJR
7kFghNvEPjmvQ9ZlDjyWEaCIjZZXTIvpVAKXqFd1ZatskJP9jbPZWg5zrnE+ua9gkk+SU3XkXStm
p1QHtW4OJmuxjCu2BJyq0fPVJwWV3dfGNVzhvd95mv1ZDiAoVFiRpy6pqJZjKm2o3rBEGYhc8OX2
tFVzdm3R3BrC03S6z4TrVlpKmOp4a2y29Bq+/g6f3EH90NV4fWLJka2aF/3hSGsdwq7rReCzeAOl
QXu5ao0rzBo+6aHSI8YDa8wzJVKKTkenG/68tOmAfVfcUEX71OpCko6T7spWLBd1RY/OSBF0niEA
P5AeWAlDQEzo9Pf1Y9k9NmwGxaG1sBU+OobCmWrGyeNrRokdijHltobvUczgGMN550N4+jOlkZG2
LJvO2veXJa/1q8ArnvjWj9hjOUfh7sF/JjxgM67CJmfGgn+olqEfiRgTegnawTnn9A3vYA1H3R0q
+hYCg74P/5yuh6gke6t5Uv4sA+ojpDOx6KhrdmKxcpxqckZfOrGrjph0iSo2Sx92iH96DtedTS8w
E6F6EDB1Oq8I4BWWROZvXTU/KS12jvONMXDA1YTfipUfUIgknLKH7ikrG9fbOQ+PLd8IjbBvjGdR
1yNd4AKlytFvloQUr0hwrr+TGiAWfDAeAbayBPU9tS6181HrJUtbQtU8hwXFbcUVGORz4G/aeMq8
X+GTjH7lDT+iSjrhR2oLUFmr+E/S4SYGGGJ+uiaYX3WZbM3H3uJq9SKLV5YHEus6+XJtU45Jlebj
NsKmvLQ+Hid+nGLt/d7JRhPOMGHcFPxJ5gH/8Zj7krOnHl3PJ9eRMaf6a496SW5v6rlVpUG8hwEw
0j2B7BsWJKFkfeKwAPmS4DXsishv7e0hyXDNBVQp/o97p2RpkBdu9lmfmROBiazcfwRyal2Jr0zf
eG5Bz9oPVHG3r9TA2Oteocx8MUaSC3o1uD5Jf63jPQ4xrYIZB1+DDEp3tEJK4ffxbsTLzglfL9F3
4Maco5PVkHK5qY2SnhZ6jZgdQzdM6eb/4n7Ix9qggIsxIVWVNHJbjxtL9mpdk+xqODpuZm0yRbou
RhC0e2oODSShm7u297CteLca9RajO71/WcICNRTX9sA5Bwca3/IJejRLAhqZ3DCHprVjOOUMStEV
RF/+ipJ0yjWZ+mdQnPgnrO8OuxUaGtSGAyAGllOozM1kasShxtLvvvSvP7Dzar3oohhOmqufxryj
eXPnfu6swsj67fRoJPgPBjDnDyc3Tww64qRYArAk2o32TvIIU2lC5ypHll3ZrkOvJCk1+ZSvDz5v
ui+dZJRinEfk8cipnW0KvGIGpDooID5PMObIlUahPYT3UNb6Dff619mWwlFl/e6TNdTaX4Bcty+F
4nozD2eb0cLtPodF95APyiQgVH+1LOVeW8WDnkjWj7MbPE9NutO+wk74q4rLfl9cjHNyIlVswcsx
GyUgpNW3SO6yhVvyUv43I5Cjz0xH+kcbHVFmcziODVZOALBtKJ2+7U9QeIOAWc7ayYgB8tSGFKck
6NL+i7lly6k3qCgyauIpyeydgCpthkLZXMZBcNUKlNadyPTSvbAiDM3TezSGinMwhozV12zLaTLh
3fVoZgkqBJnBdc6uyUCBI9Fba9AaQ7NLmKYCduAS0oCYRzCn0+8IJdc9F405YrS7xBMgwO9TxwKg
serspJVNK1zzZEmxhqib18jp+Hw4Y2JHxjw96TuGU7K/OsGi7shdGSSIOqUACPQTipmQI2tyz9Lk
z5cb66l9b3dQjbdxaNs4XU0iqyHsRoLYUUQVZFgRC+WjAfZh2n3dCKkmndrBelO0WUQxJ03gZGNj
ge2ggrNNUVrnVV9HY4TNCuNI4gpnKt3ARiJlfKC+TGxlZG3coQA3JEkULdYMujBFmkhPNwEkCJJ7
PhFJzk67RHWT8WFoKe3Cqd/JrQCnlPST0Zg3aZRiDqnpOJKROZViIMoK78hwOlKeyb/eIC97s+ks
GkHqdhneJJy+3xZ5OsefP3Lxi1Z3XTiFBIgueZzy8T2sGBSivQliwhUkwYHf37OEpabst9IsnaQM
k9Pkx0Zlrct5Nwb8ceS4RuZtC8Pod4dDD3a6M/9Rrxe5slNsQtBgvZEQyut2DGzu9vwSQm4fpp8y
C1AKePngrYSLhCfobKO5TvvLBDvdXv4dvZCl8iHwqG9NvEZTnkdKZYNNJZU2KN3P5YkQwIhetyV5
NsuMXlWBojlameRHEJvll6B5Ef9fBsVRZncD9atvbL5gTlMwbVKWvzI6TkSfDkAqGZTzhS6KpFrd
RwRa+jSlC1YgUjtEiqYuoCLrILZwSa2JotfXGJ7jCYjrUENFswgqY2tctDbIP6eRFwSV2jHN2a12
jC1FQ3iPHGNxrWcDpxgrdQEzVphrVh2wvMCQ88v2Awu60h836hzMsLvoZPikjCDJzrC/m7nWUuXV
DL8hBKfSIx3D4QTcnuYsz7UtXezPCYNY2PynDUblZv/0s1nihK2qXDWWEGTchtwIGN+V6iQF2sGo
rleY3oKdV/alT+IPV3cozOoQpB1I+RiGEVRUhIMwgEvrwEJEO0F78TlI9moqR/2JTwHjvcGQ8AOH
ZEws2UTbDCmJNyFF+/7WzDIQg06cnye/IUpCwlfZBTi0AZG1Ut2N+robg0h7BLOa+G4P+EPB3jqh
zNUnwekEyffczH2taxWm07rAb3OzWrZG/bORSqWRKmCjVKUNMkPAvh77FcUKgynbR+GC8MR57WAm
xVoAXOCLNqASkfHnA9qC6mHVBUUsXalzNqf5+CLpaEBoeNrytUl6OF+lQ0UIj62ZchehrRum4OSB
nN0VocxFu8qm+0sW07yI/hJaKegQnno4ff7+mL8Zao7klTWuh+j5Oz2d6Jm9UA92QuJC5MgNO7PG
sIGOerfqgIOqj+o339sTml1DFlh4ZRD7S0SHyyRCOseNi6SvTGn/bNjy6Ep0iyZi8G0zcOial5S/
lV0PbkIiZDCmKtmk9m+sPPJhgBrwRJ5qPhNTDvn1TMod3MihOBDLKh88FlHqX39+ACJP1SemJRRC
T2MI0r/MK3POKUC9YsETde5iXk1CJ65eXSqxI6z1qBYHMfuq0HrCoube21kJBRVdYxkD9T3+BuzJ
Q96i40N6I4IvfOLp2CK6YgxfjoZMFmOD6enqculvPLShMNHTpSv636exIBreOD2Ha9o0OQmYMi59
BXOnsI4okn8wC3zU1laNSKkcStFxNzS4xSmQKnEe2/eQEHgYew1LqS5TEEx2xezwh/SafL8jLppf
ZNMDa668NufxTsDV6+FDXSYHyltaVcI6kPQ9ySlM91Ps63wRYy7krthhZXFCV7ztBWFJmeWcTtgt
Iv+HHPrJUt4kg6vH5FvPuwFaaArXcb4CtsxZcrfocSwqbIwCEbLnjYaDSuUVTs+sD8i1PbaI4/x7
vUAtr3gdbMkX3OUpSJT/iwOpdvZYTfqhhaOYNSdk8G7gIMQ6BTKWgOStXPfxP+5ZHFiL1fz2AQE0
YwjL4mYLe6u3Q4MHH1P84aQRPKd4wlGmIfNS+Rq08/4sphaOS9idwxpDAYdgU24kl9rBHrq5pXH0
AYJRe+D9hHHIztpMSI1sShWdci6OnmVkDCGC7911hBojXrjX4wzx4yP4sDt20KzluCp4vRMUWfdh
xlnWXPOTBAWL6Fiybl/wzgqJVFLCu/PlxGR9ZzNj8mM7XbAJIsixTTUquakHmzAWH8yi0kvMc6On
mk+OG61B7PTQoj22s8wg41d7mG79O5MfH0nWA8cBC6jk0ux3iDQHAXejbTy82yhphljIJHpI9SHq
S5g0mQQ6qHETYJrFuOnRkhflC7GDPLlBLRGS/ItF93Eb0/nSTTVIL2y+z/SBiMOsbY705jVqeYHI
Ilj+Y9KkK3IVdUzQPlu+LZ8EvjqZodio1ejD+HKikBoE58y8D+OO4VOLRhk6TsSBzIK3sGK1uPoO
I5VppBcRFzm1ebZXWCz33joF/q8mrtxIZ1nhR6eppbSkXDvR4ZrraX65ZR/wqs4JPOUJXiTAYlnS
qXXyH7L3kUMChEF2nUhzqox0kWE9LlZKOGyNYey2SwdNkrP67mGEYAmMUaIGciQdgZrM5WRPueJ3
VK05Vnza7u/zgPtpEM9RgI7INVCtWQHELZpD4bWMf52RUHO4Lj8hO5R6Xb2jVp/o/m9FlBMQ0mt1
0eBb75SH9dyy2n4dXKAXAgQnRmoc4afK+F/DryWpQBSumP+NTkEob1QUTKqPMD3wiDxbyYFO/a8m
sJkqiosjXvBHpFgceyPQBkiEmg3YPilFI2fmqB3LMk3JIz0Gk32vhkXc8OyOn8P4XebFHqcjWuk1
fXIvtd0/jpwEvYMoNIT3rlOolTSElWqbnuvPf3aNUv8DIqjzCvRNvIF9ris14kdsoWzyiVCVfDwT
mGaSUXR05lfCblzgcKm+mNS/rHJT8mq7HGWIqlTVYRB3crdMgHuqclP/ARghEEJFzbDdTELWDmYM
Wm26cx+RrpZmY5lSvZtapNPLymWmhkJEg03EhCnw1boMwnP7nHHZyK3CXLKtYDItqOrItlvhmXOP
zH+cT0DLnOQatO2XsqUdvxP5e+dQSnJG59fHteaBzgt2bk1bgmMUw6OEd8znicBukwPpS+c6EBWq
nSroO6nVzJ7hGPZZkmKnJpimr46NiqShJFzAlcMNhqsUtZk/Pvutm7Hy9AssG5luXd6/MXlTjXTr
s8fxtotUdAXWOfx08Kz7dR8SKqZQPboTmRfIvWoZvxqvOYFl6mYAMtbO7tNDuJX5XITrVDG8/5ey
wmznPywgSnXR8i28M3AWcwH3fTeTzXkdph30uo7YRxt1/UwZLc/VXWQtfehZXNfo5kPiNiU7Fnka
ELMFvQ1K4dOvJjrYR7hPtdKempccBlSc8IrROldM3Ny/NerSU4TQuuMRV5xKNNprbUF/nxALb5l8
DLw2yNSUxC4dPmpc40DSIbvoAvp9UrwoJgs0QGa8lxS8DSKaTNvIgo065nB/DHl5F3IAksaRTZjd
gx+7ysqneDFhiFutXzYNY58fjxKtr6LEBitA8h3222qqBBUY4ZFQl/zLlnlDj2ZAo90F+i4K7X1b
IQRBFwtE7u4oL8cwJoFAeG0IBww2GoHA4JpyKhegxGFauk473OiavILiL5ck2OMMaEuUexCdFCMA
U1kTgp1Fr3U1Hh725hYkBWHuM37dlkLj9o2hVFXBB/77byQnefUJghyogrWsD5oKF29gVc1kDTmU
bLMb8EXKA0VEVm62Bf+h8CGoWU2ojvIhg7SE3D36+931cYeXvNL10MgkUXW8FJ5RDgu1xESqrK+J
g/t/OquJuIT18JKRAQvqbIIAXd27bI4qArq7BeD07Wu64CJJGiTprPCVPA/XnkDmvJZ+a3J96W7M
0uyur81ITwlTeLYDJcY/3RYI1fzp7lSqRaA9gmVtAayX1eyRlS47Om895jVuhzSdztnbzoLdl40R
BAiMQVVU35GAitxhunDFrprFzpLMOBJM2LGfiIVZrZPyvig+eexAxYwqu9ag4ARCEMjhLasnPn5J
QdDG6JMtdEq4ykbM8qztzx4jGecCfSccn4n8Kmtd6M6CZ4LI6xNvBOZCgqBiGzTBA+JWZwDB5bbx
YF0NfXlcWDm8STjz11XGnDsMOyknFEB+ZfsLxuJzBBhmAa3O3TFN2XyS4L531U+xFkKfOMVMBKVF
7TEdWW+peh9ToSzRcauKKdGFsaYFY4EzTCTBCuMIfHRl8Pr3R72NF/SxrYBhyotjF6Ga84xGkmQu
aa1elIXdGxeQ9xqwB75Zz8l9dMcqWVqAGriEkv8Yzw4vflw2uXTONEtyDxivmbd3e22/oKqzO4py
mFFnCRD7chmKYipbtm1Tk5wZnkl0adBX3haPFVjwo8+PUPYg60PUTHafq8dBuZiXHQY9sa0FR9oO
I3QpJcOcXtFFLndtXMdZH0xSMUD20nXMGY+iUTxjb+vBBud8z39jxce9q0TCr+GkarV96ATyATB8
w4afr2rVaSbijZc8vL3ii3oBl/jwbwn5iRcMRW7gltKOxPFYE48wVZXiye48Y+N2kjM71U6Z/g4s
y0L882GkCAE15SzlcRlayxR+S9bq0nY710jIoVBiZ2H0sYAPegWMC+Y2xHKGnIrJPiFmpvPf2px4
rLzC+glY5y0Ylqcnr8QUbxLtUSYWCly08qy4mtbFM2FqUx5+KiDSwrtDIpwBaO2IiA7UsE6UVhmS
LR3C2BgQXuobGRZLzyowr07BcTZF/ePT8HGhynEQotTZ1ofSLZcLiGwd2bSYWS0tKXzu/LoPoHGg
9ieINLIYcdzYLElZOCI91I1O9MXxOCg4qr/Xh6x6rXXTHXSlt6i6AGGwD/inGMYvaUtfKVzVi4lB
FLUiB1itlzJFxD8VFasdzzMXHrJaMRV6KNuu73r01zC3w9tIawCmHs5KOl8iKW3ZRws6YiG99xJG
3IQYN9VO7TyxP/GqHE3qjkEcyFFImuG7UWZ9Q/lCwUggEo5ClLfiKEAgLN3aL+n7AlNPU+ejftUl
PLw/CdWZbFB/noPiqyYDfbjkUSONvzP0zYDVX+gwXidwqYwHca/htstuxzRJvrvkCwIYV4xYjjcQ
aDHfACnOJ7FXvY8DfAXWeekxprZ/BRVOsbSKVPQf93h53vPaIpWnY38W8JtwYyJSrhhkfhVsapbQ
6ZxxqL583go6Mxr1BTS4LbQfZBPPGuR3c9ywT8FE+QK2YV1lp9TwPF43Iwrh8pWbu8sFYAJ0goou
fbRyid4d0Gt5+sTbp4jZEbgrmOThUn+lKMe5+7D4Dda41aMYj2pmWBoWJcWg7v6xIQBCzV2Zr0gO
fpbJJfRSt9wvW1AWjjDqmiNORMEzi0rxNeIxSz5kbnerIqJz65bTN9d7qLRP7VVRvih2Zyoj4Jpy
iBu6Ln0twiNVOsF/+GuPH4zdU/g8Jo3kqDZcjsKEUeo7oHCgzGd31KPirKy82yRgOcfDlHHWP8KK
gRM8iq7WD4JH7wDIN3nBkwf4WVXfKwaMQ1LmfjnY+Y6V45BRRc0zaIoSGEcVr3d+CTmoSVC54e+G
DXMxqSuAQuJEQPqzjzEFHkJ5Ciqa7Tss6FSf4ULadOZdojUJNc8jzCmT8vvqN6LzI2bjZtQoLUj9
IgV0ilSbFwfAzGUDHyFh4WzF9QK5Ajtke594tALVoJ4Q7BytQIb7oK7XT+7L5p/Y0z+vVnxk9gvW
ZAIA3Exxwqr2jtGv0835v9yvuDfYbWPhcJxw8lYUlYXtFYQbtf3fgDTMoO8ch47uL9iltr16PMhu
wkVY9aibzHxvSSbPRQHVBi6uzFdFo45mn2IQsNAE0AUQZVmG8iRylBl12llN/aOzB7t2CvXI6Ovy
DIWcw67jv+UQ/nUJW/Ce07Z4ebFKYr619SHfmIn7qY2jprpooxGnW6/ZHy23GMFpt70hF+RcoFFf
APpGy1sbAtEZDJ7Kd8AFJFusYqyuG1nZx7I7Pso2ezr8UyyYHPHvvliD2//dkIKgx2Rb7aUblKyT
AuRcwJVLB/lMZHe4l6DU2OayvupDP1T4Il3yz1TL8C0bISeWcUk2/i9mPBoU5V9+HFKXhE2XNfEq
2oxPS2Oe4kEbyylHNtk3kfr59K+68L4gcSu5G3YmMvvMlabgNq9O2NmugN2jN9KYYfesu0FJnRLI
LoCQgzy/eISTaQTsZBNgW/8YoRM8lkyfKQ8MemgIkUPIE6ons/LL1F/3f+/CN9bL89PHuuOSTxjl
mmM680LXspMMExQmVs0lDuJWXSveKKytltdvJ8vyMsOSgSnpEvZIwuvIkkj1d4oyxsDqjx4bQQdG
WowLunyZnRNBgWWlk+Pt3B6Rl3bchjrb5Sg9pIL1aii1Cpv+HhA2trvNLzc0YaT7RVWw53iRpwVu
3lEOnd5VQ9NyamFlS9jB80zv8hOELdmEpH8i/ArgOlqHdjvnNf7BHXtf9U/uEXAfU52PIyxaB2sH
aId4I58uPC3FR9y3wzycaluPGeIkHu5F/XF/ERGiYRU1fOzmFB22dovUS5JaM/dvrME1c4OUQErp
0zuYYmjQP8vxnuB2JmHVQnDYOM3Fi3ZvGMlQFBxxPnQ37qua0rIYWj5m5LhIaRSx1OhKqu1sLkGb
qerymn0kC7s7A8hunqKw+pfNJfIl/mgbPP2Kg1qnSD6D3P+4m5g9tzR21GIgtcv8qz68lq04q6lZ
ecQha5agPgGfejMABb/pBTJZ8KZxVyUgKrnmy6SXS263CMWHcsTwC2lt5T2zlWXGd6pIIiOG2l9N
QxyM/UcedRxRnQNpDUuHS/7n9TMMkWtrpwQY464hUeee6HS0ihdcBgcSPw99VlJmzg3nMytFz1FF
czZ6oISFvKajUP/iUPoZ9YnJjB7W/DGdE6+omfHo5Tx/9dXlJfvWZQpmXUWY5aflMFdbbfbBXawx
k+u7l+BepYMRCcCmWnsYXNnKGE+iQLZIV4iLq/dYVmpfF3FDbl4RR6KjDpENTMcER/B8UdRQdR6X
u3NpAHDNMM1m8GW4lmv5N0hu+IvsDJijJkJcerU2X4sZfRoWX+OeLrZFJy9TRMZ3Vx6rpHa25DHu
vJfFPiTTwAhl4eiM2TrDcyNG2C11vQ/igIGGBB9y5TKRYbfxAJxGX4ZGVX+O4LzHEc6EMSHSTax+
Zgog8xfd3qtRIeGkfdQDcqY0Yo4d6HV1iKPfmSjk66SJv2CNEfJaB7DoEWXstwkUEgqGnNAElJU4
zFC1WPUjshOt3yIfaIYWtMSEqJVNc9oofoDE4AoTRSEKZKYYQRoDZy5YlRk2xZbvlVk1VyR34cPI
0ga2muiFIVcRS5y2QiY+Jw+dPm2urG6rqWJJohYAI3o0rL0lAN6nwwFmglsdum6gePZwGNViu9Nl
NNI+lXw7o2pxeRtpy2wWcGFuR9GsKLmYgDajrwu3EWv10f/G3ECgcTNchshs48HntnPebhtd26+c
TQPR3huXrR2rFZJjmXO4JzA4+EBOyaU9S5SSlhkspiKlcTHzBKfTFEZd3Yd50EfbkWEXw3Ei5eCF
9zfmWG8rNFNMgnTtZcfSYUj9afIsy1ZRFG2awzRjRqsXESS+dlRg9FS3vSctU8913rycvaJn2zx6
TZ++MfE4+WUoN5s3FtPvB0QFTkE8vu55kG/WGFuwYS2DHD1Rl2jykikGUz0e/ohPf8TWntX2v4ON
9Cdb1p5yZs0RQzJEpTHlBHZydXI6iT/gBa0EvS/HhwoVCo5jz7xFi6eJ9uAcsJflutH67Fa1l/yr
wwxi9hH1b7O5oON7hPQVM0CqYcGNLZ8jWmjgBWhT5p/1EabRvc5qB+gQysPz9iS78+REPzPek+rZ
zyMxMM1atPMAxHRXF667+2CDj8Bd8+LBObY15vLdJkQbdLXwNY++hMlFhRF6gfJwKJGClgNs1WGG
cN2nRW87D0AbDWTHPe/NE4THk7NWp/L440kcMW6HOYyaGX17jLLNCzt7hnbMw7K573UWBnv9f1IE
sOEWzBP0ZVV38OkU0UqW1frx3s1RH8qTKSocapCbase0m3Lbxart3uoY4TC+zvwt1SOOOVret1Su
cMJ7M2DVX1LrgdR1PVOwAg8xoftlYxeVMn0+NJeEHkY5gW0UTiwJTJixnZS/BEg5QfTDDBE0QRAF
L2gYSpIo8QU4SgbEmDiF3/iUmbF2v+UPd1VL9F4CA48qKPsEADpp/el2EKyC/wq4yrdEAJky6jAn
TODSDvFR8CLvaqN8Vbg+zuDrTgWVQP7DJ49vMpCq0BkseOW/j9vgCFaWoQiCqnQObnNtJb4cyDmn
XNkngMvX21OsYWeWwo7Ow+bJBff7uqAAKCDFcBBjhc4YfH7uXUQ/Kb21Kso8jmXoeFUIWtxIoHlz
3z3j9IruzWL50f0eKvHQ/HjybNUoO3WSvmjX36NXebezZW00HERE/pt+DjXBIwnMtyAZmft4/J/q
grU2zG4S4XsNbnVdIHHX1vMUQxyu+8r4jtVOTvJBTgbWvDAZTB5K63m4NchmlMhjP9jiZQkwWwRc
1MPQt2wR8YUyp/of/2nJ+UBWNn0c4hlkdWyF3DUDIdgsrQJVfADoyjWe3ceZLruaHchciTk6F2wm
oOIKdaCtwfgbS+jy1eJ87RrRl6RSA57vjhOx2iubPo6soZcRt3L1XF6ghvrzxv+h3Dq/dfZMedbP
ViRoQ+fxVqxAYUBwNrb/6NdvuWNg178lBqnpxdp2Dfq5S3Dwh3cTT7oRt7l102GIDLzvS+VqJ0m3
CHtj6usUji8ianWzDH3wIaTsIz68jbnyQEnIJ0WldCWt0VJ7DP4GJ9og7yFbLrtosnvgp/dCfTx6
dQ2zDSny+hF6IZNW2JtzxSsHxo6qd8ymw391cFFM+1MX5HleXbmBkRqN5fx+Fa+LNzaNIEQ8nDjJ
adLQ9QCvvIjLsQ4B7j6hE9CqmOAJmt3JCuuP3kkAsFfI65B3Nun0A6kaXbFSsU3O3nPWzIwKw370
TdKc+YyEI27VZPszwtMapo26wwcy3Rs/4UOCpwoP/WzCawMWU/zxp1dN0UuY3M/cMFt08r6DeuJF
QJbSZ3pcLAV1MB7KMjMWtsiAfsSLIjW//duDFR+Nrww81DKseMu53g1vlLBgJ/SX33/kqw6dDHPC
qEHlfnQbgupRf0xzx+WNBIFVddbXUQavbiAZxm+9/Uk4GVXERFfyU8SjyTz/FqUjppRbPtieZ82I
dvSrhRlN1bm1tDkGbMz9E8jaAUn6SpIO2HxyeXx+R9Rb/oUT+SchKkC7/amxlQQ1mRTqHzCi1Ds/
aXGCXDYQV1TV6LhVahpgGFU8BQdo3/MZeVPHGnasX/nos1j7dyHOc+H3nZKEqpklnEYQqPLSTSWG
OSc/7vpjQ2ICe271VpZ5IOXdgKwPP1U9XztHVv01rHC/LULTJkvV3EXm/4qcgs8+mApcXo8PvFk/
9jsUxhrqLug57q3eTqxxOQ/TQEDMnTaHkLCoNqMyFPY6JPIR2agtl6fon4obMfeX3ZxDlBxTB3UG
OKpIiwfUcmhSqjB1+RD8gT4mIn9j4Bv2sXf6tMzsN9IRZyO73kX/xvTIJzeVE17LuwFkrdBSzc67
OTkhTnZetneN9evDOITZwYYGur4RypYSKFkY7tm90vfr73rAoQmaRIRb9ELnhnJWLThamtSWaKEZ
vmfVMbnw4BCgTfa6L5jyAWbUTRfMqxyJAAqEp5jDQ0btFJETnoXsqNhoASdsacNJO311DvTlnIQU
tNeRPwEzfwtKTYJKmb8voT9oQlOtX2V1RhLBYdo0YueFzX0smilkfGAYOvGoP0zCO6e5rGCeIPFw
kiAO3N8WIoflNwaN8QL0wV1662T+lW7tQuVvCeJA0OTU/0trE6QyNDmq+2RX25TPfSZtRjdcuQn/
0dNYJYZjXd821qmfRlBO4dPbfy80LtKkwm+3H2TfssrNU8EiEn7DIlPmAXqsfc43jbPWkGgjX2Ie
xni4Lf1ujNU9HZMCrkIZ+eqPPckA5bjI2B3RkKX2JsvVFivDcP5u+k3QHvma3fF47i+wLqEVHGbB
pJq52H/K2oHEQqdbhDW6U15y3axZ4ybKWut0hR/u3y8a/RhJClY3EsR1mFB1IJHb/vGi2I2Phy+U
ZDKHdt4QIe5s6ojvhYxR8EXzWpHCxHQJ7VTuvIXNWsfWGdIVWt27LKeodCBwUnkZkV+Usuv1TeBm
tnq1zAi96Giq++zXwEDGVK8T0ybZ8wSYrQHx7cAAkMfpUDUhas53V/s5ZpZOi8W9qi/iwKlKl2ZY
tFCMRgvyx+2OBAe2Y11dWHXP6CsYIilmxN4IL1L4umguzvrhiu/5HXnyj8M6x4BeE7qpna9Si4Ji
d5CsTL25nYue5+BAUHf32GjcIkaeLZfGaBl8t2UXx4MvHWg5BqRQ0oeivOrXsEXxcQxlDGWp5rRj
fViRu2LD7QI0m14NT7wwP5l6rLJQWFS+a0P2H6RrROrtR6fknCCTFxKMY76GoCwMRTBfSXNaJ5vf
GAlHmybpGKpJL7SZfQR1hLpSXP1T0n6i69VAPywUXRHcrIOnbJlDu1yuLV1HiCfR9V7lT5trZcV8
c723EYo/7MgsbXzgVNXEcil9TVaeEZioool2KM52/SXinn/WzZD8GyNW8V+5LlXiIh27Dak/uZmI
ySDCl4LUCJVRD1yVUdHlySvBeKF++igVT0dXaZuZAxzF3Z4ZqRSf4gBlQ4JBLCy7NI7Q+ogKw2sS
WQ0bmtTXCQRWnQMeBopm1s0bS9o861S2HQzM3bj1YxMzXQcKmzN5jZIGXtOcA34eegeFcxmb4bjb
OhWF+AKn9vGXPg8dQzfBiByyB4ro3FpaOdMfcsGAb3YVTT30yhNvYBjNVpnr9Fx9cuE+FVSHDMft
09AS8GiIFKA2xGKLNuND1o4px/cep02Pgj/Snx90VmtefnCKS8GsV2xvDnQQlsF/U3UP5bT+ex2/
RD1I9t9vZAtrhC5yO2oP1RaJCWa3IDSad5SLuD9LJXMlwuOwWQM0QZhgVYr3MEUNG/OJS3qmsZra
PwTxxZovtW6w3u912gxG6iNQVPlNVJWD6PCNvF4x6E8N7k3rcZkTBciG7z7FXtEQAe60bZpl0W0I
NpsVSdWVGL5CEPwk/RPDxbPIWBmIx+F0naf7bHlkH062mb9dcj+atyrGxNVfFPQ/enEPrCEqCltJ
aEQuRkp0t/14qK4NU2bJ/+V14iOoitOxpSyHBaqKlZNs0Baqypv9KI28ZWATmUbwvrI/wzGbF4/D
NqqirHPg+UCkx+dLaxLKu2fLptxVHSK7GIduMsDRYNzduDatowmqssN5gnvjJNx9EgnYaJfqPwqg
vfKbt07+ceG642QolpHgoCePSy+tddQ3P1NuLi+Cc5+G8F7c3keKsKhohiVM53vYL0ULwhUkY/wu
Dil5EfJnBxWn1jyDXwJQN4B1FRQn9VA53aYZAZFDLs7xycoj8WiYLyp0rjaC3FGVKaW31WUciIW6
v95onnh0gnhfDmuDbRU7mB523jhtZOOAGHjmbKD2JPaSMDOlXiU8ggFp4Jj6r+KF3XaialfAnEnh
Nj8zLAmEhsN1hX9oxE00LGt5SGWqN2wdioFqJsrliqSp59E/ryHMU5qfeZMTo4nFNirD7G5bmQ4z
g3g4/3VFIFUjfxgWDSCMX2DlTDT3YjEuCaZIDGJQ0us+OTpqLJrzOivvgcNJQyiuM8Nd5t5IaLK3
Frye192W3ZcdfRzQJ/lWi+v4Gug1NJTJwQ6ZSN7p/q7g7Owq+MC79nEV7kiHRZi0/z/hpw0rLvFF
kU+UjQPxlXbNpkjGZiC2kBNs4BcNJOLpcAtl0VyYdRWqlJRjkRNmNtTAkUUtiMTz0kOJHwV+JPMd
fll2X2TfnEI9V6nV+UpP068AeWbEjiNYE6HlJBRE7TK2PQLWj9iDrrF3Sphql71uWI7akr8iNq6H
/fAPiKH+FtQxV4Y+HF243X3hr5V4Phk2cJXGelqT4aIHMrBefp6W6cBIczbTyHoO0hrYFEs9glgY
cLvhY3Fz7e5TNXqeHUESa0W5/HxJkA5BQAUU4C0O1K1WUusVV4YdH5MyCw0j+XUQuwWfIxWn/6RV
BzkyNZCciD+70jKo0mHmljlbWEHU7GGhQTLR9u51Nm5QuWgZ2izioBatOZcD8I992KWoJ4EZQG30
Sl6Bao94ltEKoZihL8whgAyf/HpfBKCpOVAEyjbVChepQ9dq0I3c+/E8poGPdwo6qAI50Q3dtwhm
wBkH2TzYl2K5H53sVGoE5y7UtsRonOkgDXUUDdPURN6RZtTqqOdvQ+6y7lQ46x5AoLqqzeF0HoPX
OCcmC/JZ0xuYDy7vsirL2/ed7DiL3Lgieztnnk5XrfXPCvluMHdwH643qLkyXmUJxS7R16c8cW3w
ufAQI+gblMEhmeGLZq173DRfAG973ela78NvgDxwPTruC9IlmYKZRxo83CKvdmPegGkODQVgzZ2U
LlfBLNE1JmJFzSfOlidWXxGKQ8TC+o7AkG1DL611fT2z9W+KPWaqQjCzj2UxNznbVZpICJGPFjZE
M7M4IUWHm1tlBy/c40Et9OGIeJe87cHyzRc90+MJmZWou5C2gdkxqZ1VmP/7baoYNdYyvtRbEL/V
pw2SALaalkS3ktl49jOdkiFHTOOLon0sO/qOxEW2r2aZntHE6qHEoiFYlnUv/Grwd/4YV1xg3PoP
BcC5NQNO+OO0oIPTD4rHZVsl6IAtw8jFK+0sjBza6TK+jfivq1L0Qq3dUMh+Fwv9ZRQw+2emS76j
fRk0hSPmGB62yaH6RoEOpN4TTT2//bRR/bYasIvcgkb7gxckLQLNZFS8fYwEsinHGod1wKbStHtN
YY0rNLryZ2ILMYxl/ukemy93sjNZHE6QTz0MuqLMPVmv0uHe+1zZFnk2MG3AO5dKQQwnxW+Yhjp9
84cbNkcyyA59bm+dIyD2UiuFcEQ579AlYB8e8+johxnydGw+gvMuAJ1mbhDNLVossoAdktf3o90x
GYTMG5RhcDWEyjK4fybaeRU/Li6LhUmDTpRMMqj3XrqzaShj08C5znlm52wu6DMdSVcyQbvnawjJ
C53sREk7hswp8/KvUKKnwVgW/7rqmZlOLIy1VrPDJEI0uvmV6RHadO6LrvNKVsc419GBoX4oA+DN
gXCb/qCkVOlyK5XPlDcLg9xOn3cK9HGP6W+dsyq+tIAHQtcH0iHE5Why92oxs3UKpNVLA25ggx/3
AKvrtaWL8tdYTE3duUQWpGSnkaXFPLTsiXbEKBr/wH2FkpEd7hCFPkhr14ToO6zdKX+rUlgJhrgC
bFIuqzJ6MfyS/o6KHCHUsUWvSd4LdBNiw2Ll56oVaV/SddYE70AcZcGZMi5Uy1/UKl6DHE5lf7Kw
3Qqh4roUOcOdnIsgnfihbzdy99gM15SzlXdLC2J6fYEreYJecXS1662gsV+tsELKz5xc5wwrRw5L
CCrImTNTYjUOtl6IEOGal7lluI6xnCAx+yOb5nTsO0j1TYgkuUZzzNoHiUj2ph7ZEmIuVzf+O/go
COhfeHKKhmzbaQvNfN1y6FfIKHpzqDPDNlGWG4dWrgtZ2aNtxmtBUyWv5pTZYPy6rb5of+9FiDKs
TmfwwXAK65S069BEXX80Icvrxta1wKXNB7a2k5B1bDZt8Q0Uku+e2+GPzr8n4HAlt0V8d29507Kl
aqHAwQYEwG13BP5/SFzpdExRGOcq1nToFbZRHJe/VjscdMfkJwXjKBXrveHpjIwaVviE1jWfH6Q2
xkdGRoDglhlI5SzdHA1hhPiqZ+7VVbYiYk1oYymEQV4363kDnzJ8UCyXB2pxbVCPb0SNAwOeG2zP
brz8vqJrW+3q0qU73kIwhX23GM3Veo0xQ/zx7N1gWOVxSJ9E3aBzp/Ofap825JyLXxPmHJwH+2N3
2UPU4ayi2mrSR5ipoV2DpuYntkR+cnBpk7wAPsc+D9iK0O/Dy6jXgA5h+bHwB2SCWPZcF6WAG4BR
8YpEdiqNeEjvNVk9ScrTGnevlVd5GtCm9F+JOzNoh8IR+aW5on/9wOiOoV4NasmUtLSnhwXv7fEE
gARjzW8L/5XTYtLwIDFm0gO8bzuLNkW7loUDoULTqvQSWe0kPn0SnPzQKQltD3GIYgmURwjiIKvN
MW93p0fvTFpfT4cW9lG/xCshur4pHX6tkV7ksheUKWUAgMSNBtvBl2Wjdx8jQ645fn2kAomwpsFm
8SLyXT/DAHgfiExaNhdgEFdxk+rfVBMqHjkKIgZdgBNRJBhWYg/opzi0+6XDEDkjqvK7wFZOs03/
ecdpXo1YQcsYI4bxdOSpv0peK4mWlch7fc9yyJcG1EcUyN7oZ2lUOt0T41mh4iZYI7INTWKDC8QN
YCOMfoOXN5ewB3qqAcJSzwGY4zsRsa8jPU4TPeMg/F5ep4ck7rnFwhs8h/shYX9w1z2oCcRBmdZf
qZBn/9+V2BCCVpqYXS8fPtGOjYvIumqNcG28zxgqiBc9AxNy0988R8OI7L4eCMGlcnrKc7N3zY+n
V7typjXzRHvAxolW7/UiV6deKUaQ0d+MLz0lEv12uVl7l+46rwjYaFHCXsJrUK/3yUZ+qXzhS39p
CNg+Ib6/gKNuki91uXN3yqPdMFSnttsTD/INXVa6K8gvhCf5OROT5YO8TRE93DX+4QPqZJtZLMld
+dqVbrjoq75RtwsH4xANcbSuuvuARFFgw64Gt4AepHU0rhcatXC0ZSmmBUY2e6lteOLyYJ/1rJJ+
IEIZhJAuRttWtxz9lyPddQVbqDheOQlCTB4s/VMmnMnLZoGqAypHJ8Wp19lL1S5S7G6kRZnalGfv
7tg4TmPXcpqoQE3/AbGl3TFT+28sK2G4k9/Tn6K3saHHChyOj0tfNfiCLDDDDUeLaRxc20bOKPVp
KeqL7THOztG/GMaJH2my1T/90W2pRwQCCxkyswdL9n0XSQkrRDwk4maAWwY8XBVc0u3UahuthwUd
vy/XtITcCDhCn13tSa7hy+Jjf9xzxjQwI01HskEt6E+KKl29/RlsJjU1F5XHmm8F+IVUlID+oiuR
1h6V+LoP5+XHuthK94dHF/yMyr/NSSDRVcHGvBVsgzza1xg/7Y+8crHxDs787OJJs91uneHwQ/ZG
BUQTdHv03//qVoTXBXA2isFQRSBa5xnHzX7iZXTdjlVtrrii0dvurCverIbxPfZJMCHVNgMr/QC/
qGRDx5tdKyiyUM3nRUXOsyiMWAQFSEDThaY7KBPKwm/EgW3bfG9QljxrX+nch2rvT4aE5k18NZUL
Mdd41yQ3DM7LNWyKHpxue0aGj6y112vVKybkrszCQTMGXaV8LtNQG/GcfO7O6KrHwuTjQ9BwDwop
yPt6HkSBjs5nbiOT+dKgdXp8aJu9sKoJ0aehDFj7HmHo2MF3c4jI1Jrk2Y9fqSk1+7ZcSdZgpuoO
i2K4JeqZPwpimM94o7lgk0B+NSRRzEY0tYMzM2RDfxqw9+O8q6XfZ7hicN2HlnOyicbd2a/kYGj5
dllhq9YYEtmkxNdUN7HTMtjTui4iqkV+3yZ2GL75JW8+o2ulCwjEmGrJqr0FPWn+saKNgtCj2jUY
1QfKx/vzJ25AdO0MkgZa+1DhYuyANtW08RkEpq+JN+I6uKUpv+HWyeLp8AmKpBkTfSH+6j45mDdD
DsarxGTBns1DUYsLvM26XfsXdbn+hQn1sH5AZ6TaNYPQPBnY2KIv/IRhhLJPc337fA7kr5wwCopV
7inBjmEbkozotRIPCAn1S0UMsCsIvkPaftrWwk9YTY//cDcBGdL6JRdO6gDJ1mTOHFU4L+LR8kWQ
DpOKqbTrBRNV3drlM1/BiOFGP5XC34i/bYR/a160oPVSQM9bbBGB17rEHWuxAXeY5BBlMnf7PC/g
i8PitHkIcF7Sm5SD8OsvVtHvAxQI+oqiHhSqzDT57F9A6Tifpuvaoco6UTwepxVZOP+lqGNR1ijA
E3DpgrOTEsMQVEeFZiKKYpM/TLBTms2Vrx3eDGHPYUpKFZfcdNKSFPO2cvHd2cmzTIjYt6H99VnO
YuvsZuZxD9gLmXO4PqUv5kvnUxBiVzlZVeqPZddzG14uDdaNLC4UmvqMrHx18AFz4cbKmfAa4SqS
54/hNZTM01Y5r19R2VWrPrQZFirOCNwxSHTUnFtIEwdBQ0qjR3RccD8DtYa6/FOIZ2TrZi+rZnlu
s767z6+wubDsCurwERy1yscWXNAb2LcqGREv5xa6IrhdGPYWh3OFDKDQv6GRRCNBgakj8N+VRFlM
7/qqSrcDEk4CIr/vkFWnLZaxraUiwk7fi22AcjltD3WYPE6c5kP0dp7j5ZYy+Rr17WoxcoBLs+0I
EyVsKE0YafLMmVUdd4kzbKHbmcMjq50BCM5iFqmVr7idGxghBtkbmMzQGROA3M46roYCH2rQHRuK
J+uTH8ZVuYcGEMgGYQdRRuAy91b+WkzOGFuTAxTygDpfaVpmxEH35GN2AzE7t2dv3EKSywo9ZgKe
D7/i2vLAQmKLBhD0P1M46WaspAmYvXRDtyMjxjXAAzFxF8isV4RDP+njoFxCfwp6iYPHjAGxya0I
Kx5QePRGOpKKUldiaQS+Fo0bjAPDsgybGPuXWrxo6VEjZAQZvFPV4EbaI/ee6lPzrIh/DVX9XbK2
6l9D+Xl4iISP2jph6O7JwdSLJawTQwB+RAGcB2qCqIvxGxvjAWDvlZF8ZBpvXN2I162pUmvmPYjG
zchwBTs/gsM9jPbpaKJSNnMs+14e4qDEJmoq7rKRfbizQR4mji77pZVaGId/+kVcdE6WrwzgplAP
RuVnB9Sz/9gXUaUtNqvMoen50qiuHPto6dwB+9qYaDHdHQcDAdd3eB8Kow+EHbmVQuVglzxGh1XR
9vdgni1rgufpAF1Z1wEIcTaucRcpB8J5VQhgQm0opfcWyAC1sF8vrhtOT4oIcYDFo95/MfM2gWsF
ocs0wRRQtYf6RDI8bNmei4VtLuyoHWOnQYTK4kLk8X/qAGlumzThVMU9ZcCVlDP27varOW8RTLYG
+NtEvy+6rM+GIGAg31DqccCbr2746e8Mf4y4DA9To9Pq8J7AwsoGNUdZLDrknXKlKEPDete9O0nq
Oqbs+MCNTIueTw7n4AIHI6WgfQJCGOZS45T/tWIUeEZuYhw220hGIgwD5mFQ9Mg9R9NtyG6gVKko
IbCJnfj+SWCgwSfyaZIB7V6UD/iuf/WiyijiBRDQ19BpZmFNjSqYbJYibJt6VrJMZh7wA7DYeFNu
9S7VHl6p6cLQE7bM1iMp28lWpzijpTQhRy+6xq5MbaNriA2WMtn0S2jnrJEQu2pcIa4pUS0vQtPe
JjLbiswh/b/6qbj9z7Gx+4eYv/snRmZgtlfFjOjQzdzddpLV+atrlcdM0BwkEfgDicpTGfAmb1fW
Z1KD6gphN1XkoBogDZ8/o6fxtu0HDHfp9OF611WNgZXiktz7bq0NfQae5iY5XJSs99xdY4y9hJBg
N9TKQ3NiRJJfZkdNYDDikh+3kKft8CE78Qn1ouiAukxchu6sZh5TAGToCNJ6Tio0H30bxvfeyLYi
SdO/hMHzejhSsjG42S+auO+8GKJP6gLcCuhjFEuJuJ932c2T4aY9CQ3ru4PC2N9x5G0P2d2vJ1Zs
8QslgdeQ4NrPtf0+MnwFNBq/QZ+rBlgFMd9cDmC5ODgLNBN2g7RhmA5y1/BUZP34CTe3jqYdJBCP
KLd4y7Vv3EtvcEPq3mzpVCMnf4b0xuJRgwZyhWieUktwF4QE56xsuugeHweN9jEXLE6//H+cJxb1
pophQEoWSGTW5Ut7Im46JyEk59PFzVRowkAcHyo5tEfxIk3ZKTrvD161aV+pGISdYyYRvrneSCnH
F7LyzFxq+ihEoQ0MBybvwSv7O1j0y73n/xqqVsAMPGzU5nyHM1pzr2H79uCdMGixXuF6bsRn1eh8
3//DgcEAHojRion741TqWkWxw3siVG9PePAyRumrMxAmSqkL2rjDd2fEk+aqVtj7pCVxPfN83Z36
7gB89dOABKT+yIhpx4Pe0mjL/hd1BmJmfbHPZqGQ8mjJrMsfbvYsdRhdi0XIEkO67jwIF8S+TIQR
nYkqBHp8x6Qd20BLsqXjWYmS/Ngk7eqNhxHue6k7XVbnN9u1pielI75p0pTc+sJXGTSYL9y75kxQ
MO4YF9yEnW630F2haHcO8/BbnUDBSbKJD21LaW2Q/Zbc4vPo8oQb3AWc1LMo9ic5aDmugqr+Ey1A
OyLJzO4FlVKlsA0ORAbI+6Jexw8Sz+39JXcbZxWb3BqNG45t2XYav6BLdx09rM+uPClPASmt4mZs
7QM8wDSHhuxbcw2a+V8BrzyajtbgogHA2P4KV16R4dAzKd1n3YBBBOi/RU20IQ0WcJaIpwUHmrIA
VCV5kGmY83xJrlZJC3vanxrKOhJr85JXb4S63hJOiIjcV16T5ZuL3qMX9luUOs8ktOhnJRGstTYr
TTr1XAsrdL/c/HoTgxzB8Jrsuj0As3LxKF6k13mqLxZphd7wDloc01OujoKnq+aqOC/Q7glRjOu1
l2B7q5aPA7SuFAong+xfrn4SZagSAVX+y2mN5dbQecnuzojvc/dv/bvIDpaZYVu/AnT1DD1V3UvQ
aC+SlsTjNQjElebw7mpd5uFR8jG8kKZ8V6LD6OxcTwShuu1kzi7l/WXveaL5K+0p25EFVOgO1qSL
QKhv72ZTO8yehpSlbRKxP5/Ec4itBztWFWV+1dX52BtW92ANXSTmrocuvLAz1DhIq1U02nv2hMFP
OjJ5kYJpb0slNN1rT142+gdNQfttHapHuOCDVVXOjr056lmE+4yE6mf+02Cc4V+C6+cIS5MTCap8
bYyIGKGw7oPppzil/rKxDJhivGWCKCkLgB0vcb/YlkoVoypGHJqVWTenqry/TSA6I63+LAUOk+d3
Py4Xh5qnsgT7dhcRpEeK0vc6oM+WfYPCZsxXScpeiW5iUhOvPztdGXKwZqfnT/qMvo2ZhYGBB4Ck
MYp9FWeLkiVgdaSTWHorevcZOCtofIQK+hv/flow+0ammB9sZNkUsgcDIPygcgUqUAq9V+Hqvgk5
/uW2UhoYgcchFpzz3nOoguZ5eU0YXd1O635POJmDxp4hKD/an4LVKLTQlMaq/Jd8G7D9Jz4U4Hec
7EFPD7Yz7DjKq+9V/ul5ia432ryCUzoZZYPxxGymkBgB7WpLIPsYt3LQZ4kKgH5pGQruvUHO/HQj
/RG41fAgMi+HVnGpRf1UfaxeC/kkq+HZotiZIvulGrxtiscRks3aBHa2d4fDWU5K03zysPrbaeCL
xNy46Zpv00asRNOKTNj7EE+15lN1DuKNydVpJzlPe0tPGMP8JSf5YoT8C+CxETM3NhOY27Z5v+yc
oielv3qc/eW94foMw0PFuO9IWz22jK4yVMDy6ACubHdu/FMbSLFHqPes1CxDwh2N/w3YVMFByx0A
Kkr+bELM+gKmjslmA0R0Sz39VmNsC791NK+t7OjfbxRUptNSNzJI24S9F//QDKNcGoOpL51DJFks
lxlFgqialyft2ZhsG8T4hKK+rmiYxkHuXNU3b0ml1aUEtvm3y1NdFgjsnYNEoSJ3Byns1IWYK3rs
qVd3ljZ6oJLxgfsYDFzdhy5/csxQmXikPhXZYDwTVFxv/Hz7nVtTD01FQ6Zr9/ObTj7den2RpWO5
xW4R5AKOseNtJfNz0QnmSWyp8I+Xfq2QoRyNoPiIyOZAjaPpeL67BxzJHccK/DB8uryweE99J2FO
4xThU9qntmVPPHgJ2+uFdkm7ZlKuYBH0691RVROH2FbYTbNrD70/2nuTpat5YW7rOR/sFiXY/K3b
WZ6Bb5LLJimJT3E3fM9NAq33A+ePPe0OX32MRi01PT90oBuvSUUFyGgNcNvRQGCEDT2ww887iIuO
FBLJRTW/AH8xvDEWrZO1uznWqVnQcWaNRlo4xZIf2QCx265q75GfoyyXTAiu2ZWuBKnY7zSU9N8q
+wf43/v9d7K+ajNR9o5y4ugTJ3nF8FvNa9CShSJ/1zN5FXCI6hbQhpWa2AmVzPZrjQgwCGul3IQ5
TXvBvrVqYwJlZ9pJ4DuaGTCG+P0F3YRP/Y+cwLMMdHu+smFa3PH/ZMZhQ7tPD8sVopF8aMGoBIMJ
++sRbVSwqHMfCkkNijxX/5R4Yn+3Ed0k7+Bp+mndE8kDYC7l20vKCEFfsZUojjNRwWxrVTmUBl1D
l8vhyeWD+ejAoYtO2ClaNfyxyHxx70zgCB+EF3URAVeZQUHkwE4xbtBRexokXhfq08G5/zGwa552
T8gtTk9vyMuf7yhXK/m6DaAsVStG1TPoScwl5uzRbjPDfnfXE/L5X1CjYHrpmoRTm7l2z8cLg2tc
UE8AbwQIlP0wrPlmgDNsCr+gDaYAbNGlHP+HOtoSRVcwAR3aWyCQmHFUrAWuGLHGUimBCci2jphX
IvaO9TYsXLjiGwc/t8LqVOPrrbOABirGxYgAZyZy6g6JY3llIET4bkZKIn8cRYGhKZnvJ4sCO4EK
jJnmo54GObmtgffDyAtp9EboeWzHkMbMNVPOP+Pb3ned4+ydPqO3+q4QV4R5qdKM6p6FS7OTX3AF
ujwo/NMgw8XMDnhr+QL45Ibm/BxLRyf0XpcY2dnWgCvKrqayCAm+ITehO6a1pequa2pGyZykw6Mr
xbf9KdJFtwtu3CxkebOKuCDQRtUhdDEm/hHFdvMivWqkjHZorIpLWbWfkQCuBVT87xxX/8NOgeJ0
JiaJXT5GTkeyL7xjQNhvFNxqOpmFnkRcbroFc0lylta6tnxwoWTk2EPjmC/fAkKfJ3gH8MP62yVT
2nGvSdxLMVuQxDmgzIvnfGHHed5Ym4ocflKMVvRHzCMRB1Ym1oSywTtCzwpFnSlYGAIBzI0WRjtM
FIIj2JmbK0NvZ7s4FDfUyxo+ngWpoo7BDHVltafxDNr2j3hfhQDYA6XvkFefUWjVk3JXX3Tp8j1l
HCnEeG3wW/1GKLrULlUYzn2b5J4A+gsnIQua9VBKXK5CMZWp8TX9oY2vHs5oCdWHtAkfA/9nwkES
gNl1BagO2uy8fjakXnmcrZ3KNqz0tnL/j5GUAAW+A2VhLbcH37LMktcCdvVtZDMYSdOoOyzljmq6
BLuerELjgukPUPDmDNVf1WxODhr6VUcH63vx/F1mgJGTsjkb5mYg77osMZUxfzvbgoNzREQDT6Fv
kj1Z8DvC6UYJ6P4zG4jIepBE+yhexvnw4QC0rIdrZVzIMsx/asXTi2OR7Img9ay0XzKYW5LzhDPV
ijzwkuZfiI+P9uc72yl8RqO24mGxMT8RhrZkUukkMPdTO448IEFLOCve4Zpdl/QgJTocL/M2MIRZ
+iIu3Fw+daPkik9gu++59sH6fLDjTkQ2pEiWyHnmGBS1qHLPif/9/FhhpzS9WH/e5qVxQ1AKZlgD
dKyRYRD++pMGKXEyibAp60RBygnchpFpx2VVTTMZrVL1o5efInJJpjojrUqidk8jdKrr3C63OpCp
2kXdVxvL4HPuWjAa05vg2cYBtsB1M5PpsZNVnXLbRQYW6jpQE498dJ36WAYt4yO2/naOyvcd17dx
KKNwla+cYAxNftJkhSBFz1R9XQcqhUs8BFuwdsYD2oyWjhrleHyyci2cazDEAFHVqant0uGPpRdA
yqwRU3SoldQj1GB8S3+Pc5QuOasFNd5++ztqJEXfwdHGrNhOf/nlOmTKNJvvqEbL+5HNRafIDeXg
vM53CH82tBXYW/xx5hTfYhzTI3pK1+vy4vCXlS0FScrPj8gsCrXCM8z7BJzkKEcbNljAdhLx9swe
Y5Wj6clAkptl8K7hd1m7RO3uInUvCF41VteFfxWHOZEC7EfD+I9P2CReypm8tkgaSriAG0XIZGqW
42To2GcOyI4MUDylTGSpkEhgroFoE/J7zXt6cnvf4e26i4XquufS753Sg7rU1zXmmJ0Y4fiKIzAu
5sJHgqTpMYABbwQ5JP0m35JZUVD5WdZcZMpSo/auozmUqVJ8GGtIrlj5HEw12o5a/e0x/QMc2vVr
QU3ww+TffxX4mZ8lNMFBRX+cKdel2FnW0EK0++mArR93UO6DTnW+8r7gaKahRIgYFkltTQUzs+VC
/W+aw4+JbdijfVB4F3dBeyDcXfbDQUeT8p7w/jPUgEnLLCweEyp6HEopsZxcVH8MeZ/wH/i7u4KK
8HBmcz6fDxiwG3sHEa9l/ad1AD5EXAfxGpHx7ZUHP8DEhfsMfBIQ1bmUr6wcbPl6YZf7lrA4pzwo
u8wU8VjzjahfY7R4D6wEBNsJdVEdzut/9DQDchNnn09c5G7fQTp57dwNX/nRGfByS+Zfn5CVyKbD
cX3E4T+1FdpSM7Jw7vhKwhoZsRxC2reGG14ZT5XuVJWQ99JGZr2v1zUFXjBwmIz+ssCZigJJ4iVR
Sw5j/RNIlP/0g8GI4Wm8fvWWek8IwaWkHcFrfwT9q4nq8Gt2CA/UaYyJBM6rzcF1WWTEjm/lOuZK
hqTrbCHnYDvrHMBr+XHKww++x+u+Z60V7whvs3bxtjLqb8VhdKsC5HWgv2z88Uvih4e5GtP8e6k7
jQSgXf+lh27jTcCE2bowX9XnGVh1UywJOg8I5OpOn2MI43z0pRZxi/YM06x+lrBUuSCeVMwBEJqO
xtixI0VBK0pC4qsWYusqs+xiC6gFgYjYQezBDo+RfIV5HBCPojLYE4KJ7hMFUTDye2ek/UgsixcV
X9xqc1ggqLbxy/SR4AZ4imTj4uCdi8XrsWu3hZxyL/CbgP1V4N4iFT/6OCEvHW/DrSNTPMY8cErN
38DwaR5tfsUhglqSrACNGdzp6dUXh7ymGRW2EXvWyi2+SIhPYMJ3u+N1WayrwtjNHf9HuPpUAxzt
sv8hYZtnfWPJT83HXPTpYokdHtu3mCbwgB2oA2bbZtfvyX6vDi4479piNsmnpuCj2q2jG4I9zmKR
MLoEzh/A/k9jQ+Y4SfSQv9EsyfYuzCylMNTBRIpBTp78n14akz447gu8DQJBH9QK6bSam6kr6VAW
8jlNmNQ2p7YTCw+6Z7lTWPm6RA6t7ZsICz/ACG3AVAc+N380r8UZh1QgBX07awTI238854TDQvVl
UuMXsekjinfTm8nbS600qP8VflBQfenByITc4jG27dhRScgUeMVu+lgQy99YrtTju8KpYStau5RO
msCZx+kq4/FmhuWQB/wOEWHWJWRWsONdlBWdpLuS5Rq8NS9lNRH9zcvIY676x6qnQmt6VdJQYGPs
tgUIUwoxaY1+Ct3qCcX8JS/7wjqer0wmn749g29QG6IxBWcjLHG/KzfZ2aKOFUD09ftM7e0ZqJcF
2My1Ln6+IXJ0xmY5vkV40KoDf5LLmH6nvlyM6t/weAGDwGLxf5CTNLe+G22GVdZrDwxr/nUk1IQI
gqPxic9T8NhJgLdJiht7Kfv3r4BHg7ZH5QCWK1u0P9BLYp1GKr1RLLbxytbThWNmJgUFSwV4gmm7
R3Lt5pEY8+D67bn/nn0pVb95wyURGZ7jN+pbAkxTUCtQZQ5eA2Jo19GIjNpi6CmaVOCDDvGEdWE1
+4Y3O7XrDJIs2W/Td9ApWiMcfzago4PAMGWWxrTQHiJithSudpBI3Mp2OPL5RV3ca2XTfs/V4Wq9
+BxyHf1CB9jYwPvFwrYwpSLMritKGJQcXD1vffpm1REFEKbKGkQ6A4FeEWfK1+OXpcgWiXkLV7b2
gOVQ17RVbiQXrQ+oDEdujbyGb1EzEmJ8XeC0fsNu9kK0WPI6R2YjCmvNLYDnV8ybNGPwH9e+nJlv
/njr/U2kd4UhAhPmDRDs5hCFAeNONE/7Ow7XXdZ5bH40GexZalcO7hNlgccIMZn5vnZKik2DyDYU
CJHNCa5ll/dkoJOgdEeotrKNmrtKlP99Zxdk1tjPGuerzpnhMq4/wNL6NRQAnEpQd4qRaeB3guRY
M9YHV37smpZmluxSH9NrwCtO6OMl3FIFqNDjp0xHhM89rsAp9AeLFT9P5xQaF8XqOrSxTkyZU21S
OZo3S+s4OThSNcYCIS76sLzw28SPepndLkSyhTJS5OTwdqhXqDLAE760gSIrYuCaXBc1DQhNAkkE
ezOpNTRPua52dc+aJ4zvA9GvnYEG9sA/+0fIJ9m52rABONP5pXeq+c5TvrzrhykGM5ey8jb6VK3P
pv6RjaOdETmYuSYAOuUsCmLA6YVjd1fcfxhKVu6DW+YpSv/zRtTPuhRWw3+5PUQ1HT54xpe1Z637
NTkmEjctR7Umm8OvCVWj4SMk2D9JKQ3K1esZmzV8+ajcH61oAYI8+KtbGGt0ys5GT4o7ZZ1lnKXj
D/4CnFG+ghxDDvYrk5cDsflUz6zQbFod+R9Zs4CGCR2eZIC03ym4K0jM9hhUvAmKUSGn1n26uODp
ESrlH1KSqZcW/FjJ9CNMnts4VKUKDZzwTE6PlwJAy9OSDtnaOoM6xjBI2sC1nX4dVNErwR03B/ol
cb3mJwwBZfOTykbtM+eEG0eoXLZ7J/r3noVgYOhZc9Wm/Xz/hLOw/GRF77p8hcHthF+/1pARfDyX
2q5JxplEype21IijjLtyS6qRHsmiFeIpOquMf1aXCzzIwkkrTb8qKRGoGROI5mG7ZmqdcNN7VMPg
O3EkqaV/slx+nS7XXGqczwgxy+Ruq15UrnoaIYpxMNd+Ob+q8kNdeFW3Bn2yWb/UZFNJDt+F9hwP
NedF8GHUy5BeGlZV7ovw2AujIXmAClEcE0jU5o5UWyMXp4Hz/DCNv2BeNuYDzXRo+7A4n/MuqU4X
rMdzArz1cCLWGZlmDWy9v+i6nZABcR8fkZbWxdfJyMXjOD7V7zdQHvLxfK3yW6D9+Rog+YER91FO
H07BXfBPrQOY9wV9k/tVr1pqd+r/38KckdKrXy9Nybmn/vDxNRoTeJdS3ZCshi9Vy8WnVwZjWrat
kjvClrImLY2SodQBqG3s0wzO+ity6ACLUGZ/dwqjR/RoDuEr+490uU0A63gZ4u9Mam4QPs0DWAkE
5hKEY1ka21Xp5dFDAbUZ+NcYhA/0/TwXkGprHsMlg9Yo91PouFxb4GYI2x9ztUSxLF+YmXE5I0ZG
xw/VjaimP/QI8tQbCm7nQoHdJ+Qj2w61QY3T/lLu8ZFs5Gby3mp1pQ2u0xHazEKpuWtvEfmgRKT4
wCvqUPUpImTXhtUxV1FrGUnFMJyHar/bS9vCEaHHesex9qbYeMxsIuM4tQflp77Ml/S1FDrnf2F5
cG42aOZMbmieuh0VsVvJxxK44rTA+mK8XTV2uTYuGJDnzi57Gt3Ezdaj+UZ1cPWDEidudUVxxrDq
Zl6fzUbZTOaHPehkPSR1llAnD6U0tem7E1FX3PuazXfV8mGqGiiW5OjwnGUqRCD9BefFqvE0f1+3
Dt3d7zRKjfKL4tgvIXHt9Z2LVLsdNZrM5Yyd/F9qzmFmgjmoCKdlUT48mYNSe1A4YOOsYAq1JTTv
VA/3lCDTINPB8JQEm+e1q+4L5MMmp08mc8JCjlm6H3x1Z0jFoagnmmjHnzn+GMrYPrLPm+5Wk1bn
bGrF/NjUZlhnv96aJikYW3V5lGxgG/c8NfUOSImlEJ8YnHgJ2bWhfKPpb0Voc+SBVeyJGoD8SfWv
qrigPIobwC7GxQe75HkRy76Q93KDnTbdMsWI2qgBu32XjM5bdu4JjcUb1ecFeVv6hFZ/lMzygqeH
d2ugNTGpeGcdq7DJ6CO22gyKo5ySL4dZnAG5bEwk0QuxIKPPGsu+8anE6ycvN+6M8bCZz+TaM5Ao
3BScAN4HOSXz1x+w3g4ELnHIu3euGJr/AVB7zOq7qb1Y6Y6mxv6d17+0VocauuPThLONKPzC12aB
4B3T4yTFuyqjfpUv6isLfruP/Meu41hwrUl+8TVrwLxfHkkGQXt6+d1+QZJ7b6xhIPWVjfSUDxd7
YhOSe5OkwY3l1hu63fQa14K5VaKaZqArM4S/B0fhPThKbWl1FNu/JaOBpi2E3yc+aZOhE+8pF5G8
4Px7TkscvkyO/Wi9eEuxe0MXjUo3quHXNoWoygIvUtnNcdKMB6K8BNZUcIQkJ+wFrLcnlAKYYzSv
f7n8zvTuuj9yu7KaQVJekOkthUm+sBt1nrfUKCYeh6ijma5FAAG3RcjmxkiM5skodBi7K0qG+Co6
1bq7ws9XwJTQUUQTCCbBod9pvBa4U8bL79XMSjdJgNgX4TJCluBJb9+PbIPm9H8Hzd3wuFRaZ3YU
j4Y/f76nyAkEDD0uHI4eDGtvtVl1gU3FKcphNpVniJwzYiMmAmb2Ht/SNdX8W/E33vlrkc6O14VQ
WhbKQ/M+Jihk0WVcG6ycCfXtV8NOyAaaHraDqAxB5NFQZWV007/akk7tS7diJnEkUYW/3MAQaYVV
6J/TJvwN0xVadOs6E2tgTXjcjnDEcvqpNHqeaKye21yeZa6SclNyNoZQ7hupXv4t5ejwoDbx21K1
wxiJTUHQLw5nQclsuqQNhEoDrzfxeiTPVJ2q8zgipYE3giEWzTMeUoa0g0xRMcMwF+CLwStiNpuu
ys+0o9+C9CZrhG9BYCYPqv36dwgvaz+TFwZ0G2KSY5wWKh+XkVkn6YF9JHoZRiQ0f5ANuzP9LRSi
uBnDj0YxAw2SmZolxIW05V2Cs7zH+peQrB9XR2+8nVIgdRRErD/jzPz6kyXXXN1PBZGmpE23q2f6
AzenscprEDbLPQNgtdnfyrciN7TdmfxETf6kz+eVjsO5OMLuJch40AvHx1ZSqpi9GR16QJnB7BsY
epNDwLxMjCUMueNabcHw+MdhSMp/iSz5tKEUCM+INfY7rnRneFhA7BM2hoApqXL42FHewoP5F3PZ
Vm0nP2D5FI/DrT0fgd05soMBgKaM6xIeu6DR7YHvDkSpyTVxzuQ4Pd4e1hjYEASdE2bw7210KH0K
NoAp508Oq2+zZanufp0O+hOIbqv/w3opc/HtDAQSNh7yAasDOqNDse20eR3mqU+1B+TjyJWlY8ll
DKPw2F89cZAD4dh4X2+nhdtKRlS2uW4F/YbfqwObQY71m3Ji+uR5Ag9NJ6emUo9DeKo4NDsf0fgc
e7v//KMdM1EaTSdrtHkxPj6qHSKN/+htNv7scG7/g21UWBzjO/IcMqJFye/abmMnI0O06hEJ7RYP
G8BMGoaA4kYVLfpdtz10QpAYBj8mWBU1auSk332QEBmSsw+lNmeYOfNlIrdHtLUbY7oMa9bWZQMB
88/tQpKhUFvr+FHd71qDMpC2PunN7oRbQtXd6PhCIVXU4iZeCIlABIySFZuvNxOPeuQzmMRkqmq1
j32tPKhnTEaOwUnCERwvT5Rxv9GwVGUkxovqzjaolhhIKcauP3n4ePtz6PA79UmC5OpOX/2yXKd5
gLqQ8jzszXXjVuu+zUy3gA1W+kCyHRA/YTuTg5vI8OnlDWxew1YPdLHaA7RlHv1j51wdU8SAw3rT
vYYyL2ybj1iBERX8nDRgYf2f5p3ciz5n/uiq0reDNBGAIL8bvc+xqSn5YggI+GRQfKFVc/9x87ll
XrBdY7OpAbI1JowBUnnYEAEebpJcw+EabjaAa9DCtv3yiRIKdb8+/9ymvFGoHgeMBdXZMe3SjgWg
+TECJ1GIMr9fCpujwHLlexvPex7LvdiSconpOJ5lFCDmAkruILDa4/jc1yZaiR7kkjLal4psfIlR
DvZeRJryrkAWLqvSvj/QymqcQ99WS9SQ5UZwSBgFCNaYVyoGG5Mz4fkRR6922nXmyBqaKciZk0yI
XJW1JG0Y5lEjLnV19vPo7cWAWZTh3xoJ/NMK2+js7ZjTVs95WIyIR/ZqAIr3wjR1hqpcVmn2Iqkc
myl1EKRYKrdZyf9efxdd5x7BuSHhlkAQ5br1Mdf5xhcNISdr2YOLYZGJQt4stCySVN/nW6G0LuOy
4f4qCdm99BTDjjQdCi1oBrU8fAOnJR71oC5YTX8pHqi/itC5rRIXT9elZj/s6CaUPNzIhDfoAgwp
U4xCR38k74N9u2ZP7ZW61b9LiNsa1h6WWQQ086PAHsaR6Fpjl+dYFFVKkKjInOAsh7NBOdBujFMS
zUGXjJLcyLKv+RrsKly7RKOHAfz63VVd5AHQrQttc2dUugphYocW7kQDI1OcVuPuOXubZoR4qZ1D
8KqbM5RN55Uw5EN29vXzBgRvR+whwjGJhRI25yKasYw0/kIx/mQ/cfSfIURKgfqzGn+0++u0VOiR
nKI1W5qCHhuJevnTGv19lss0KZHSKi2DRNwSGhUS171XAZ+aOUuGMdNfxT/AyiLZTOpAqbOtxlxX
i8SvDu4LhNclc9ahLcgphiaLZmK/GS8Jp+1OpWTBwSgHFwze9CRDrqmhkQ7EN7ucHCT7+6fJKb6r
N2y2V1rl6W5ybA6ly2atwCiCMdmXiyRT7v9FqEHSLPg8FUg7VQeVNYCtPiJ7C6QR6D/+rJkhv+Ka
4v7iRdzglvwBj2V0uUbYUKZrTS5uinMZnW5kq3s0cfPMjrrl5WXqaGPUxet+iFBqUtP9JhFVkNsf
DhE9tGsQ9tsyA7TguNRKg7VC6okWtZylAAsI3K1x5Jw457kulE7AKsCZ/hcOfBWSYQWE1yq8nQly
8beQa9RjvL4o/CdOsCfBQRCnPBAb9o1ziMff3i31jNmFiP1g/KBmTNf+opV+tRRWgFLWVV0dk0BG
kio66ivD+jWkOtILWLX9BTBlW4MI/UUtZaxAlWEyFQKVg9WuVmTBq/mV9xroHormQFKF4NF6o50y
klGKr3xZNurwMDhBMV5ccFEUdajLvskn1MStP6JXOVj5akypyq5lMv85Rp8PDjGMkvJa1Ki76QkS
VXfbkdjHu23xSQGUhaIjBPUybhAaBBN0jSZFA4T7r0PO6rZiMBKu1yD+IOtc/yN9kL0EECM4wz0X
6Re6yEJSp/5MoSkHiS9YU7xtrHhtwO29wCOOyiqItSemQynmXQpWANE0GW2mmg0nesuGH+YSjy8W
XtKaajf3piT+XxeHWA4pLVwr0AufY212bWO8NlaJjZ88/luifUpgYMjymUN7r4dmvuCxrcbk9l3M
7xJZvXzsf9UF1aAnCd2o43sgYA88okwYGhSrtKPYGTPsXyytKt3EuZYWGUupmu64IS5FZiKOPESk
vTni8AgsP2bGbyYrUV2s5SJj1LdXnfgu6mMWfiZcEGYfGA5fyWIN1wc+PGT1viTRQhyLQli6avyP
zv4NVxG3a+X3QtvqEK/tBnhr/Q/Eu2X1OaC36gk0gHA5QMIZIN32WLLMX+v35lBoEcCP7tsLnBZ8
HHbFsXpdMVOadNa3K+TEHLX/TjO/M1pEPR2ehwShloHoqftyNk3hZafOS+JPphZohBtaa5nNJrBv
n0hg5gPk0s+7piND/bconLHAFCqVMiFwWcQV9fhtoy8AO6H6QFQUEO8fr9UkaD9g/D+ZZ8WOFBCA
zyD6GsvMkdSHPwMsPhqmqwg8/hl/slD3MHToDXYSD0bHSakyWd9Ue3tkYPQOyzS1gcIyRT8/b7K6
qgO4ujgvy8rX24WoOnBlB5nx4aNRRxSBMyPE0QjIYttd8XSFBTvyauX6prhbj0YQOU4GBNduoBdf
6Xtn07mIugH0KiwFXj0h9JlYFaBn105OkgECSOasctG7BC9H1IbfKw1oCAU+7OaVn5bLBU7PvSiO
gyTva1lihbMZz5i3gJhKSpww80QYXcfBgBgnuu9Bkv+dvBUfYFTEHZPkLD8shCHVd7sDiHdMW6zO
8o99PocJ3rppnQdXLHJCIAbTpaXybyF8zwgU8Udb1n85O+ztYqjtTYEqNvNuBCMg3/wX4JM6rq0l
hkE4qEDXvo2TPgkd68Kgu4XGAdtHypyyKXGDjcB18j1gUBvw17VYcEAQKs4Ogv7EZ9tb6nN43Vz6
lEqb7O1mWve6Tnh4dJuyjbMXSUcSOQmFOIwaKlIsAtGKZabbg39KG0TCqeAsNIC78juCvHLASnFt
c7NTYL6wXUIary8+hE/wf4adyyLeBMEk+RB/xI4hwbOdq+tNRDf2XYjxbf45q6dGMyOR6vrrrs6+
Z5tXBHvDBAuk3VzuFaGPl17kNzGKrexi+Z/NC+P6iffIEyXeEzqy91yI13PHARJUK24iZpMPc2EM
nqCDVxGiCRFSzjkd2uxpR8Q2IQ/LgYxwiS+ok5TpxVDYf54ejKoluMsFsOrOoPcwW/vl2B0/t15w
jWl1xxvguRXBtvOYvLmi0GcMfejMIKSPX9COupgrmDrzXZVrymFDuDRMSmCTf434/A3oD184ZY3Y
vzssgLldYHPIeCsIkXEIX7VPiuMw1IaXgaGzPbdl8aPzlzCieGCAzuwfA6eO4O/h0YbTFmBWq4hz
xlUSmEMS0yswrcxaiO3P+TchJyoSNGLKmoG/lSgDmxsvKvGNznP9IFSURwqka3isGhNb9MIna8Yd
gfGIXAECWdhnOdAZy1hIkJVq4qDTx3ho6RA07kxr+oda4zTui99/UDpRTe+CRMIWC5UT55A4p2k7
MnUIsKDachEXSaffqVbbhXWDBO3sC6oERAMRW39rtwcUeiMYvXz0ADIcEjlyrzwDebfhA1v9GJkI
/mmBark8Q/jNGZZpTpciTxlSbFq5vBYiVmgTSWBDv3Js/gvLOGXW8AJ6hVj04xitVLqeSPuqDGoG
h0Uzc6X8U5OVqSvtq5erMTwmCbglXcWIQRo/1KC7kz8mbG7mQP9aE4VRd+urMwUro9TL726dCOdR
FPpHAagzaRGpjPL/AjS/hknD3lSByzhC6BV9f9juQO4xBQ0nqiLR4OAsOZ5XmwfqDFhyx/nlNtML
x3MUloPowC04fnRgyXiqSwCQBEJljsg0fB34Y72LDRd8XNzAdHLuSl5Szbxz8P4D87fR0EyBnY37
p1tUmqpLmkMBkCrjSIghDRMmtaNHxGqbYAtx8Ekv1MzRXiclu2Q/b/Ebpv8g7Cze79mTti2/7Qpi
Ar62335K5Hdk34AR8CrSvfcYAGu5mPV2x7YyC3zqeKTEnsRUB16enLEzcKttsvaDlP58ljTODXK3
FA4pRX7MsJ5aEQClQ3LD2b765cVHvmDuRfDc3RfOGYXWpwC0O3QDjPw2AFz+Y16W/mx09NCrJ3cw
fAiSjD1IG1iAx7ajaQ+sL0pnVfNwkvsoq9pFhhvZ4JRyEMkN/0KoHPTO1yrDWTzWeWTb0Cj911Mr
o7ps0rWyZ0OULkAsM25Y/3GPzbo1agocI45A0vh+jm/w0qrCfWH6Baoq3rR49EDyUwlHkv6Riwyg
0QkMQH1v6MoatFSZB9SLPTCZkzxWdYiVnfM9Izw5OMtoe3IWY45FH1R4ZYq4IRdutJBeZtRI1B9e
BFE9q4YDRSr81cs992GJ8PTbZ51nqq9mUj7AtF9D/193Hanjge5Pa/JftrNA1QQB75Vxylw6T5RP
NyZoJOO5DTODilJTOHK9aGpXdVwDBJyz8MKLdKht52LGBEB82r8I6tfbC/FhND2zOVlnBjXMJjzZ
D8GOY0YzTrsf+8NgIAu5o/dSoKE/FpzBmVN6FpATAHfjex1lNLYPIbxaxLI+XFg/QlZO2PW3B5yV
26/f7GI0aU3BeidIeD+oVfskiFV/oQZ2UFgTYxn1zv9r+swYAJ2uzk/jQOPDLqTWVGxdqByNl4iX
Ftp/D+TTWzON+gmxkNu1SHFaetODp5pVopjtd7JqGS6waU/1rhtWB1v1tdJjrnFWE7WS7PC36pNC
Dv3CP+iWRVsthYrWJQpupdjIkuX3rzEUvR0WQOZHZGP06yb3X0f27ERHM2VAATrUxsiJ9cDosmAI
Pcafg9lfZzxvydyG3NUTl8MRhuTfX4eXnXZFvo+vzIO0rGhRjFxmS7SgcU+gmasRctPEr9iW9VT5
gSbsB27c66rRc7CaXh0kddTwSIxe4/S8qvosikD3/Bo77idrjY/wWMosnrd3aX/iDuL2UZ6IlY0V
ClfeyzkLcIkQrwDB1gioLctAgOeBWB8gx6mhvMbyIxgO9hi9QN6vlYFSjD3RJJxGEBbh70is6DR6
iHR2lK3JJoYJz6UKW82CzvSU8MdudmBQvzvx3o5cxmxk6r+OCnlj+ySzeduJaVZ69r6PJ7QPTVW3
fY0BUPjdG0QipB2PVQhZhhaopNh1lLT5dmK2uqU1UVDZO/U8poyLFKkpX/IOeI48P7uo7KsrXPWC
XFthyYtCqoSRfUnZIuHtyo1Ie9g6fAWGkdXyGxr4+640o+vgsnDjOEf8u1dtR9gGryfpFPiLk0f8
vJ7iHxgIZSd6Oo838+6EQ+nD7iCE5j/FytoKQRleFOgyCBkGUqKHDuZPlxrgcXjY+icaBiHd6SpL
HUPryeF8WcN+kuw0AFCvlMWfUms7b4fIDNjdrn6a+u5wGmYVgrV3UbR7Y+yCajN2hibh6vOrCmvh
aTN0pFZjHywncbebZllrp6qc7W3UB1Z1eBCmNY0umGe8++RzUzjZIH3tpRiR2a1yqVfgqep1n9DA
OSCBe2iDKN8npdv6mtQtXT/2vD/NtOSSzVTfXCoNY01L3P9ZwFItmZBM0M5+d2ADIbFWR55FC6n6
dRGpLXThPWD2NSp3Hbo6bWx60OH9fAL3bp3p0fsvNz+0erQwuOPCM2zAxzeydn3tagcBsx52PICh
XjUfeoqoNfLvnjlRLk7aKGqeh7FSuOBeTNpEtFixV5ZjgMaMv0jfj3NuFK0WrCkSA1wqlbKUY6cL
qp8mBYL42HC4lApTTCrqEL2hsKFrGVH0HdNy6tPLcgkonU1cAm5OMyX9afeIb2Ij0rUW2ZydJDzS
gHrW7OjsqRF2HazrEWu3yChapGijdCug2iMov6iP6UhJ26m1POBzPI3sUWQ0maf0rNtOsNrkqZxN
EsIGsYnd4ZQk0nzAME12hHfRfDKsgs1hDtfERmqYtUOV83x0w0szOdft8X65mVGPykS5EE3ScRjQ
9YY05XhlV6ncdPhhZ97Hevv6nrnmD/KEQrCqG5k8g4/47LVuB509KrtWVDkNNS8rkiVA8anqXF9m
0LLwQu5/GNjXOY+ENEtBc5b0pfXxZN/TKGYXAJjiZClowgbCuccv1FVnur1CB4ewE4BswFsTVGZJ
W9GZfol1rEhKyKoZdAA4n1oRbngmcRKZM4ncv0Vst3YG9RfhNjwqkoJWzgSezk7Mxp2UkYXJNMp5
Bn0ibr9Uxj7MzgBwObFq0OR+rSav9y9BBLTfisfrcIrqj1Rs5FrbHuijhsqow9D8PSYinMiutiUC
GaPtNdjfwu0ZORKT7O+e+bmIPiVoBpJ6YHRo341bEpHz8mD8uR8MP0/HlEmVwIvRIb+utADUcd8g
DR0VSNxeEhXR+chGE6tTAIj08W7/azq7mxIoKzNJag+Vy+xkhzB8F4gN3lj1DXaopOGGQB9lj4fZ
b5aqZXr7Ti9exxf0P3LNIoCp3j6+6fb2RWyOVGr9v346oaSqxQ1c6/BnDY/CVee5fSL4PKzSE5VR
RkolXq7EW1cYOneouYG9HkNvmDJr18dpXumttox5a6f/YDh4gg6I/wIVTSSNrQjkUNgHSBzaRKuL
nwhOVJEqR2pNBrxrjJPdpTkyDrr65uI6AU0OlJQnKOLwp7hPvLpvqQChue60XTaWUE+RCpSDpnVY
m8GMR0zetMcigsqUuapuOOdfRdU/s7Y+UBL/tMYiMriS4yNSrezbRKjm92kcLnnrwfovale5VnuX
iNDA5ziZb3gNGEck4BmDsm/Lkn7TphvoxJF5dsSPkPzYwTz1o1Ar8xqIxctkeS3Cggr3EJ5zfJn9
nf72p4O/XldAj+N4aMhQd+Yg8bHt8U/5+XgZzwsYFjbdA2Zb3Tg4J5Ffb30SaUsS0YbD75olUvV0
0Cdp5Hq3eiVOSBSZ8V49Gqtb83sPozPVlaM/UFvsz7rXLETPcqGHeR1yljn5moE8rI3iIDcHIZw0
ZiSlpPwvQ7kcIN7rPAvYyQh6ut9evEPEkmpr5vUm4NOMYhbwD6eFNzd4TJeovcUdeNvdRql6ur4j
naem5eKIdwlFgW7L9jit15doKBP42afi6NLi44JNTTlF7Qi0PyoknCNkzb9q7/0I/XASjYCq8H0z
M+/ZMSC0Yo9ldZuWinfoXbHoBsaDNZiseyHxIOSNSe8aSQNpJBr9ZhC7dzJAPth5kLdPqf10ct1b
11a9VpBKwq5Nlqqp2qW4dAu6UzKpXY1EiVMXHFDqqlUazfX8A37GgtE0gDEum4KQLAKu+9WtRl2d
XTTFC8MgenJB1trMZPXUc80203nwVkbRSppW7s5+eEDB1ftIWJBbEsQyZTQHUFZqMj64asUqcs5q
7BtgngIEDQp/YoXX/EOHjB0mBF/LLUvjVUVOft5sngfntSFwxsWEGxLuTFEEpGPp3qbN0iR6GVdH
cZSLyky+/gxCdH7ILYkbSLK3XPfTXOkdS7KBqISsVwifV+dytO9637eoSa2J2T7WvcdD0MB8lSCc
u1pamKEeNS4BAXGuTPJko+RbjMPbX1sD79DKlBSzuqE26bO9r5G+hw75QeoXkPvFXBHVE3iWdjqR
if8npPYkZVfpl7Jqnl1L6XY3NumWPeEe2u1GFBWVAxSGJjBVKukFSbkUuxjkiqBhMeJ0R/N8Mpda
p6wY8q06c67YLqkFGRFBX1rg5ziIZQiI2GhD9T0OxlIxKPCkTlAXGHCeCFHEFfAY2e+rGDdocibI
qEsN5GuihS+vmhO5dBD9bzgWUlAG0efT+ENhG9REXG4+uMlUMj7D3IKvArCzMYigzYfROHyX0XZq
wJ7pJVDadBVPr3KwMOd+6VmUEvQanV2rRmYNLqba8lM3q5IFbqDlzriRgVz3NuPN/t2qwdyB1FA8
EShyav+YDm5RZMFAyPki0fvoFxrrD7wjqXzZzuICdj1rlo0Urjl57hoKo19hSXd3eqp6ZR8mPd7c
UcJIaPh3AomI6IMVHrHV5GMjh2pNVvtYUilkMu+d559XAKdWwChoieaS3lp/Ddj9ICaF/JDqndIe
TabIsQj3yeEgGxpth+AqmrtWyfpZzhhuxqpk2ZVXaQGuzw3za4Juk7CkZ0agRESq0bswzfiq+0l1
Cv6f67E9wamM55bPmlcFDeUE5yxyq9UhTqT6WHZw8u9RM74vYaXAZIs+ApjCWjojXBfRYzzyGNaN
T/bRfboqpw4IB0igbzabrmyGW80NPUEOOo2yzyyVjOoqhmVQ6T+fyyZdn6MhvwWh3yFhsA026Hds
gT/6X+kciClRlfFsiGQBi1XlFly6Pjsid/7PRhkVCHsTgSoNKyvM9tLuJSx1P1yNxBks4m36J6g5
CzXIfyYmQRGTsd5e5t3osiNe6F49gDpl3qX/ZQPVFg33FW2BB6ifxIT62eomIxT5+oSx86cdJX7u
DUuSNCIYv+rRwElPetEzag23xOOyrSYl+4dBImANamB3IsFykMC8vLTxpTFxQ76SnB/5BgaIHAQp
mdULge3+YUSOXxPggSBTCCGWzGkj2KgsiFSjDUZ3l8dtPIWOkWcCjS6qPcvtFNltgQ2zLBLRahJN
TOWr5RWgoUrvBWjoiIDRYK1GFJRaIeaMS+3AmAukvw4inV+glJj1AnDx5fTdf4IroF9BRIlr6OAf
CPLRkzBhZbDkU6II6ssWppC6vDzP7ZedCtu3F17Nbn6btIn6bT9rEZhRSkFcjn9jLjBRjrQG/dWl
2nMgnhFbOvsoBQne2Aok5gcXx5RoLkUAGyK1R+fQjRgTwk9oMeXo02rqpbbA6LvS+l33GMYiUfUL
uOUABMlz5jdKop2Az6F5L3O/5UxhLnnsuwc1pyAyc5ohJiQ3arwT8RNSMSdSyxK0C52sgEa0WRZK
JLH+Hg3eMdBynar0fufW0nRrxdm05leV/xFKHgVh04mtcE02k3I/eMGyNR5WECuzXOlauIFu9eka
ekENJ3dfEW8+3S0l+v/8Gucd3EuH1Oton4K7LL4Flb3zDqLfL17bLr68J2oIRfYBvOX2WerGNYIr
eRoGZSP0BPL/zdL/dsQKeuxdRTSROQuTlzwrCeqEZUBYK45XrOGqXd9JN8W8NQ3IzMDjsjD6hkOc
yXr1wCK8HQq+P1E473r9VQeivJ30nS6jaxo+OWaKmRSkCG6sJU7hqJUznctceviGVf2gJsRery68
inBn2Tv8mPZ9mI+2GZRiTw4+eq060c5Yq/Io1JBGb6KfAYie7dpKbTu4+YqQXunCfnnICFXss5Xp
+DtNuNNMps6i+MUvd/YI5z4z4Xx3Y7wROYrbff3QaO80CRkBWXIvKnFgUX3CazKmzV1/n7uCL4pi
0P8uuzJ0eLuZQnifTjabCg521Uw1JGEe57yYNJhvWv3TlOYIfrbqOVtwfNwZiiUfiPDGLi7cyYL6
+hHoLTD6gcyAbWTAVt/4uSc92gT/UYbhOXpbU1QaHeE4Zj30IfjkR1WyejeJdtt8bxpc78BgQgXf
eSLDD3lHNdtX1oc7hXskDM/c6ZtsZbkKBagO0zvl4G7PapQrSpvpv4p54e0422bKZlSrcx7vJPIZ
q73AYjp/idBOuQ3eeE4bWJ1ur2nXDSkZnJou0blZdf7b8C5fF1KArut9qFGxhVr6EYTxfHVC6vKw
fEWfjYTNnBUrrhS1CkW+M3DxkN+uRiQMSjycVCVVJGs5GCuZVWkiCd7xpsM27J468Uffat42qhcs
vPjmPDG+lKKsYxZmR/YMChDmRPHc4aU6eJAK/xHF364z1qqKyGLfxNDNpN9g9Raq+2Db04tvoacx
F8BJ4ZodiDhyC8D2sdrXL0+U/igcN3cN7owKXddkfr9b7DHnZbaa7QYNjvcFFNd3k1055nWKYwmG
YMSxv/RBPym9djOKilG7vBx8bCmMyXCps6m3Ins4/pbmxe2bo6u8CCKdaGuEa4akX+eseNNq2sBB
CCnr6FmZ7mO0ICEi//YsVZODIJebiw2yGPL0HHQqfKE2nZndA+KxvXDCf8BrCUoKjiAH/WgWYKk1
wbW/tUsYdf5L66WRVOvNpMQypZ1uGBXaKPp6b0MZvQPsHGxtRmpnvbYFyqFSnCd4keNhs4OZRDQf
1i5GAm1EvRzt14fE+HDTZMHsb3q27MrlTGm+oZOCFxXQXvgXujpbaRpMFxM1ocRiAjyxMQMFZ/b2
EU2aLA7g4sm0k7E3klr9xKRAZN8KhxG7kWmvxVDi5J0UzfL9DGB1hsOkDSNZ2jePJxfxVC5c+DNM
V8bRs922P2ZGjaC2S6DB3msEROHi/s19rTlNOFB0LNJ5HECb/4nulATRDtOBC8mBHFSxn95JvmoQ
oGoO6FjBU/IJCSHuaxkCeN7c1QR0MAIgEVAGGnBavakq6sgFAP9BjZxb9fyzLd9keD66QnZM5eR3
rIx5TkMW7Qj34XIeqIqd2+N6/5mWrNfjAF4Ec5Z5lP1nRwSDfvLB8kqbiv9bT9uUIsJuBUGAufXN
I7Ji0W+7fm2WyWiW/2pvVdH+O5giyPrnOvuRWO5DvTi9nJUde28UA/C4BbkqJoyJ9/gFawmkLBz/
01de0vT8wx0gd6/TsWzs6yTCzyMQ12OgnBHqqOBMQkUfbTRk7U4KYlVpJmTqn1XP9Q/vKjPivJUK
oFH9zXkBeeAqRqTb4ga4SQvDV3a5we58ctKxWRQyedok66fooCqSv5VTT2lRWdRzRHNh97nRSU7e
eEbweFYO3au79fkZJQqvgYYY2cU3Tw2amcUt+UCnyJ8W9lqYg5kJwQcGW+q+3GOowQp+2VSsfaul
I3WkpEYKg+Uas1VFJ4JW0gGBzjX7v/eHALMmnObQ82xpkoAAhPS/edvGEYBgNceRX96joH1xq02b
y4Jm/lhDtzP5nYPbCaFVHJaGgm7ijScxuXF3N2oJyzcTgI/U62ZpAQFD0xfOy7Tw1e6jQr082IwD
aYzju3Phf6ufBr9o0tI/z0OYLmjTiT0/P+sUl5jRyqikxBbtbx4LolmR2pxXzBzc392wJiBYsJ1Y
08krK0guMHUvrNH+fftsaEKgAhm/tea800qAHOlo1C82/oDeMF4R9f61aYgfTh4rpvmIQsQVmhLc
HsClVzLPOvNqDMsezo861NoTSUzLAhPcaF4pbsp1qNjbGIRUD2jrix1U389OmEGxiqWYBHXJY0Lf
iF/8a4KVRC7TVWpEPTLCqAdS9Y1J84/zvC7kxAbBbmSfoflxxPoLDIkcQ//gTV7hljIjypbHTK+6
Ilahas4gyFN6Q7SiIzcI/fPkYAePOQdY8HZcm2WDTN/8IRh2fIZGbi0AT15txI0cYCHRy4xkBb4o
zD0mIU+9gopriCXHA3O2UO/bVnudqkZmAy+2oQocrQNOSnes7/Oe3X95gNewHdIwZpRjSR606Kip
35yZg9txqAvrVH33d4VbwHHr2iIp+i7sUTJEosC2ik5Oka40yQ8/W58aEjWw5Dqpx8OHPTlELUuy
3gaOFHAcbpXEvRfb17n0aeWOu2yl4WoVN4hdw9edkZaaWO8X7vfPJFt07zmnVtFwdORcbuzOIv9E
umjXBEWG3INCqysPLwZvbL8hoJt9GqhfnUREmNqGp0MLuiYkZaxyf9ww7gytxmsgWIGvUOKbsa1c
2+oWdzFmwfamuVTDaf4N9vKIxOEXnmiuJ+zWNCd7YR+/1Sg8jHU1NzizZwjrwo5jDbarTHjYGQGL
HPAmJawHR67Keq/rwdmfrq1SSI7WFOiyi+Cr57e7tAZpz1xwmyZtGBj3617QgIWtj4ZbYsSTvWVT
sMgKaao6gqcmetSLO0H1VoY/nPh3TThf4TuZe3pWXy6THvMDTlQm/FOcfKApPg1h6YzsuWnpUJ+3
c/t4OrOtQWIvPiHbEQMsS3ImWRnQsXTl28bkCAVI+e58/Di/Ax2ry9Coz6C8sbHaF+nqM56+zUN/
W3RYNnKRMfs5LoBChOXXkMe9o11OLR3BEueD1T7r9QrfL5Im7Cg2FpCVHojlKjfrZ6cs5XoKPiKi
sp/hS06UX5Do7BVBpHq1XBti2iojfc9EjX8DBbKPQVzGXBBfKbpYECRrImyHON73ZJ8ADMyGxgZd
4H9ofPQ2WY3N08FZVTM3azDKN7+YQUT5i3HxrZIRmG4Dru/1j+AnLlV1SsleOw9rsbq8pEMpq5hZ
TNctgnm+aEaoxNTVX932BOgcSbUeHrYSVHQtDVVzDs0e6ngrCO8bMZJsFDINXt1aaC34QwZmqzsV
joCmwjbEURPnccYs7nCViphKjy9sCA1R0a5yUdB+mdxrDcC1naGS7ckPbV6Vq6b7nXApJpJ6IPCA
5X1sljjtukHB88PZD8TtVQckhsDZ70f6WmCnoG6sWAms0mYhObjyYthEl4vGLEeDcNuCxUNGfsVv
pNq0/tHFdNwWU6aSCmawJJePwPXFeJ+CGgBn9qqn7dWRUBg7CbRU2RHWMm7AVtb4mp7LChk4C5JA
OmQy+4yeyd8l+1YY2x3mBgpNj8j0IVjohE8peOR6kGrWqeHq+B/qnSn5EeCZtH6TeOHiTHCk9HwV
CP0iSJPtG8JewCRyg9AugL9PtOvhZvD0oyMRdPMQ9IiCAYBxh0+PurQF/G6F8l56kqZ6eHJE8XET
vx6gRLo86SiM6YQruOkRUC412gy8bcUMWqg3JqlDqZxSJo5h37+lrOzIo6jy6IH4oTe563jKKN9p
KO5IH37VEYF5sQMWgtkSf2vskr55imH1SmQvsTkrqKEAy5bFr0R6Gjt+yztHVoc2/O81qRRIQItr
e1/dmI/PfKyjLNv5LyjoCPy4yReqz1zLnpCIKwcJdl3o5fK9eC30zFfNVZihgeWgeKQ/zOQTrH3t
GikHIB8CNWUbg98FJDXqFIdPw0tAwovVc+hmOg8cpd7ZCvcMpW86CYpj/CwYcEnZtsArYrRjlMvh
h1pA8pJicergGhEFmdo2Q4XyGVf5mxuuX3d+x7yuSg/9hewdgLYNH9NcRwz+46rDfOO0YWl2K9LE
CUAH8NV2arEG0pIbQ1mIfZKl6RZPsfn/roRQVAOYgGXJ6tJ7bWuv0ktTb5Rcv44zq4bMH6hVDGVM
bCG2531mIuN3oFCRN0dyZGl+0dzbSBXE/qYEaWPUJkhQJ4zuJ0Wmu54RmC7GhUYNRfbpCsy7LMxe
hA7Q3trbylip+rvHLzmHr4WiO4kBIfaMdvGiTua9cLncBDxSgstrdV+cVA1YH9+yquhxswgRjUzV
KJME9e+Ah4Aj0B6pWN3YCXwRL4xT+vRbk8Y/UVc7yuyQcOLLs8V6rgzjIL/xz8Qq8Aq4We8vnHVp
SW+cYL42yBvSN5tbOVJsfnKCAXYYjMqKv3FXoU1aLZTd2L5b3CVk8uxCbLyufu6btHnnsN8obmyT
a8Z9W7MkIkSydhSMakmBJztO0IDtXcbzwB/JM182dNIH7S/5lctCU793R6hICyaNKj7Yq+Iv9X3M
qF02N9xeXO2AKW5wKHkjevNoP1ezn8FmwfwO9lBiDE+7mRUM6WIYuG1i9fSGG36MkDF6EsfGXjMq
I3u5nNKCJDhKfm2URbRO/FHEecZoTjK8XUtO9lUBi07sDJ49h6usmcGbnD9mWYXSlGnlcOhWiYAB
sKgwZNimsymQiDcrLsefYlcpKp+3zSKZZ3CaPIk2vnVKaHtOMLFYPjfVe6SUJCSOKeMpETtuhG4M
tVSxMYOujvntdEWZPj2/NYeErqIMLym2MKvUaExIP8GeOszfFErQc1lwWQ0XB5L3Vf1xaHKGNDfN
8HSDFQshiIAqhF90L8M1UptHO29VqaSatkeB9fI2QsJ2pUUq9WsJtrormj3bTdXDEJ1ir7wUhfl9
64PAHdRcNa75nbal8O+QhRsuBN45ncVXCIP8OTXPR8idJqgOdl9JjsiDREgpZJ8Qv8JG8OJSFWKQ
agTbTxA12bgJV3X7jlTSIUKXlxhYyerNAJC/nkrRg+ZT7oQp3L2UlYovYWk3/pEVvur/gZOQRMsv
o5QwGYAGKzWW7gF5vO4kaF14fIt8CBm75L8ZER0WV5J3SkzlYaTisZbwumjAQSErz/DoOXuDhK5c
vcXk8tuf7h3/gY5IGih1C8B7yRQZ/ynLTag73YeZCaLb/qqiU76jYgUGdr8HDHjpUYy0higK00TW
NJTelPCLRYrfSdO7aZDxrJC+dpBnlIsS3OxYNVJgHI2jYpPbtcRA5ZGH1J+FobPEDnxK0ruB0SXg
j/ML5xIxK5Ed18H22aydrLQo9JNEX3mvVulPG6A7qq9a9vWpOy/GecujhoZTRTcxGy9yvtgFiKUq
AHuRqN3xPdIaX9PKnM8Oxp3PiQAVUJC8bH2OZkHM0TRqn3NDUHtQ1QAX4ihcbo0RtIvXQ719Ynbw
yt1O0IfA3nqCmhNxn0UvDrPWghoUnXCWhxBv4GFnvhPvVhxMkSOw8XqPkSXn8UOk9i0aWK2Ukd/m
knR0ECRXnb0f/VjzgmvX9jjnbGeswd9ZoSnJ09Y448K50DSeqO17JfbdcFInHDGm7TKnVfKbGtR0
A3aOHCXu+CjVK/KhdCxV16tE0pgi6cnwgbRu2h5+rIFxaT3yrATqBNmj1dknN9Ib4jSbglB/9qou
m2skSo9TM2Q07OeMZxILdHQfYYFl4yR2FagFWSXGAOzpqq4LHigMrKScpOIRUfkZmhDUtOO50XlL
yqE3YzIQaCQtk5J1+sXJktJcf0qT26VtzD7JPAXuYAR5YceqEygsJO9NGsZMIfe5dkHV0/CW8Eia
9Yrga+WYHAlCbSLwVqpnACF8mbJQ6NJuaMWE9PpJg+EAFmgXOMNA1o2rFB+IUCd04TAiwkrkxqW8
YQTQtl6/XX8y2z3QHje3sKKx8scCATfxHQ23YFFx3djFBubbDDEFdqoj1St6UH/bHbXNiLTSfATg
Vr8a68c5pX5y5sujSvO7e1KK8+8o1XP0j2YKWGRy//sGE0blV22Sf/uOSYKD6MJeLDSSpQHmFTz8
CiyGEg75XGPORXqU54Uz9PObO6pBy9Tw/emTYUw3vhIk5X/oz3to7f+j2hBZHEJGOiYl69cCajtR
XtyqFbicyb5PWjerWYK+QgEP0iAxJVMFFxcUmFSdz0BqS1R8GVmUVk/VozYgOYn6UPX3qen0NdCz
GRgFElnaACKQx0b2CimcnTIJmOg9lXfja3RGrL/6KcJ7bPH43ReNpqbwNTBJx4TErpeOFWb/8Apa
3Px7imesXdvIDidQz5ENerqqlcikapyvNaKV0/Uf3snHfgLhIoXbfM1hpIB6O9xZ4vRUe8I5ju9q
Zc4gihbmypIiPBe6/IP/PeZiBpIhbNvN9a/H+dOl9LcnELTZKzFvI8fKnBrOuZE9wD9Thm+IqtSc
M+WAb76DvtJG+FDiWI2PA4aeva2mJZc8FfZmb+8m0Pub8aDAyhrY/CY6+OqupchfFl5YiufqXkzH
Hra44u2xt8L5hBQJmEhLgoV/3t1wFge3qVNQfVMdnXT0i1qfKO1tr97H3B3zh3BT/OsOL/Ha492i
d+z28wEe0iUMFJIO3n/gYyBLOTZ6Jtm1oeHuXTPws9+8N5nrw9Tonb2sXOXoLZiK2LLoeO0tNjLh
dJrGhJqFedQhtD8MZKwiwLodq0S+sAl8j0Vlxb/FL0aWVh6x3oeV3dBns8opVX0ZfF9TIYmWTdwa
rOL7YRFEa1mDvHHb0LCklhzI0hFHddczg1w1ir/c0yfmU/8fsK56VbGh260P2nFrDeTnFqoRsiLI
lwF5I+yS8GCvQEZU74wxDcbOCqYjtX90QbyajIDog4qes8BT+zbF8Rp/p+sx5f0nbTQflePAcAVd
zpXcx375VrhF0O4e6UeXnl6jLtl+omLZqoU0wAIkhqwGD+ySz7jvAWUP/YFSGIJQrfyVOArLWBAJ
28A87OJbJL1YsX+g7CEPZFuEkC5C0wA9qKx1IuIPKOSw44LSY4JtLImSLrJ4BmGVIs8PLx1gYKJO
I8kAiD/yg+mLhVkgfeM7fpywhbDoj6czNNUbMypVrO3We2CWRiZaQ7To/FgZrGU/LnPVTtcUXfcD
hFr38ScgD0TO+v8tYcw4/o2jcdEYeua/mKNDEv8B7BczaY6f9QYebeDOb5P/blzYCc37BP++wta0
npXd9MXXC8BjCbvZh1P5fLk1WnA555NYFs7So1MwXeBIbdBMeCajocSE4lk3Mc9YyoJ485h9LPHO
2Rox05mnoowkufbUcegyvjeGL2zT5S5M3pgAk/kePp4MgYHB+cqYKX3lxb3umCh3Ynm16LwrQTcy
mWG3PKzTA7/nqWc7othSqz84QGfOqpDX/QITmiPTyHOtlt9tkKlG4ntewV+Hlt9wk3RTTauaFIs6
KXfVzydggtIqYI0NjNYR+bFZzgAAVs2hymi1NfVmE3Ptcjl3u+wmdLjswXBbqJn2TZG3MUoKOyc5
eoHMzTvzoO7N0CSIYmu79ECFBTjxad/RugeTOZgGg8liOzZJbxgdPvh7c4atsCiHriI8dwBNA8r7
at5o3Eq5Lz/j2ZuQnNF05b6LOKOl+niMTAjkYoEI5HDJZLkPzFEAAeQvzGdzfh+3cS7/PP/S5XY+
kwYAf5gbhr8RZYRuI/42/jl0tHHBNH9e5uHoqs/7V+J5mzeKm9MjD0PYYsuP5WUJJXhon3HLyTHy
n0xL3AtUwPLreSW5gYej+vxihrjmQuZdw6thzjvPzyc7cWQ7/tnFAB2azkWfwxHtx/AajmLCBkJl
rwyMBWgggaAcVkWJVBICxjk+1/D7j2YV4Xdzh5w9tANNdc05t+EW/U4G5LxsBvj3IDxn5oe9H2XN
+dge/pTvzlx+EK3xWiZiyChp2AIhtkrZJVmAjt2KEnJseNna7XDGovepzWT5TiQbmUI287r4Tad9
uR//iGeddlW3sa7njK/iemTWiMJKD6RGfA5S9MY3G4Mnn0YotPcIve+Mmzr38t+8U/7XEtLzLxa1
zXb+GGKpwJzkFLDrFWSQvQv6CDfLXsn90tR+QPUniCoXXBco/2qUqGS4mEDL9EvCLNI5VP+Rboqd
AzEPRtuIxEO87QKv23/RE+8Zq2gr1sCeLvJAdanztyRGU1D6IGSrJg9q3JiZA2KDW6d7nJc4UwjM
meJvJj4ooEcj9jcAFC6pG02SRMsZFXoyvDxYB99BDUgkcwa8jMebiSNwc9RrBLQpvSal0wlg+SAI
qmgGcWBKOd+ptBA/KRKIaXiLl1zglhj0JNRgFHLdCsSiiyvZnsHJZqcVjgIf19MAbAHXVE8cTRTX
N/fKzfdUj2uVV0GOXUJvQmKnJF88qTjnkRDCYXEWXhQhvnqWwUdUKVS3vDT5bhIH1J/9pcYd77fi
M5LAoZbtVJBdTQSSiTuqfs6TNiq1NO8jDdzr99VO8PXUiJXte2r2hV2h9LdQTSWYzC3UYPLtnl1/
V4VGgs0eK2X2pmFE84DeOAcsKmK8YkVhiT4vK0Fd6AGuXGEXnHjQFbsrjFcLAZH5I/iNpWeD+Y4L
If77DrNC4GP4uTlg9JIgWLtAl8O7ffP2ETKRqub3j3FX4yflATSXTDgqmYkcN8zKOVrtLsDdPWs/
cB8x718/B6fA8NB39VevYn357cbv9CUJK83jtfRzhJWMIK5y8fHn2G7VlZqkFONh2C3bkfgV70Sd
TbIiyqgWIvenKhrcWhzfPocKHVqKFfeuQaNaX79dlGiQwqxyGSEQQwl3X5vhAOMtdaKLfUsJPzIi
J8bDCa4n1xBgN4DOLWLzEb0a41EMP69IH14Et4cSBPSs0SULpfEkom8zrhN+kRZReB+elsK1DQ8I
gODcmZlLwIfAr9Md8seKkn+kPNCFbYjLjkPL082ylwjmSXUW/V0tT3O7RX2znfogN1WVgCkBuCn4
nfCRg1ldsbSbwW1pldpP888Qqtz0ZBkgA0WeWWTJoxTVfA6L/lPA3P2WJHef7D7fqfYgVkDkyPTg
hV2V0avHs/SSPzw0OLi524iGHBc5SsxcsMuE+d2VESUdqwB4clwl/uSfE78WhLOHdGaV09ClTv7d
dIRx0kunGJztvgOqcZLZDhENGLvq3rkNOIOviP9spUMIcIXbdQSl7SRFHqmnwicCU04AG34fCVDC
tE7gWbmHME7pBaXFlUskOc28Dm0KRwKaoeiqGYGUggW3bYnvZ9KKjBCl8NnxUqKXU7emZS+eTPh5
3K9W7hmU6Uya17NWD65ftjiyDn6wwF0nlKZEJB6ULz9iGC/hjTJkLTWYqowBoUm91hAP3O72D/hF
Zea7fTljaM7Izkc742Pre3urQLaikOwUZmFaaVCIh4ts8iFdImHRH7TEcwcqmJeNFfC+qcVOlKGk
FeDw0XKfmeZZdudCjtmO2o3YmzZCATekvoGIDKcOETIe1XuBUqU/KPFus2RsPQwkVlRTNnEIJWoE
w8JLLBhidDBs3NQ/4fScXh7LBfyffIborDUaZfuY6IEccnDnGy/xFjbqyxUniVmi0lG18Xb3Ms7k
1XXBqzLOhkB0gIyEyVXrDxJBN7g6VES+9AA364ljJqtd9CeAeaqO38NMQLorNae/RBPouzJWPN6A
CUVkd5I8yr8A14S8aqkfryT8wWhxLzG3KP0D4UiNlSJMsGVgs6eLJTaSWlfKkRgbR5GW1/J22cFj
6GHbmAGm/WgyiODhDuisoICFubOARK7idPw/5jUOuPX1ggIscslrwFf6B8r/FxOnen7QExilJ1i/
+p6wj0n70b/rxFnCYFz8NiI530GCxyN4Ups2U+GzSYn8/YKr1Lptbi6Uw23tzXaOAWPc1I7dEkiZ
4NlzsFIhH/EhN4qfb2n9bYDObDYs8un23HL2h2ks8u2ej+kK+7qKLBVt2VOqmAyHKGM7WgEsWlQ/
CJrciemWVQEW1MJAKJWrHyHpfWNjC6wJWksMjKjORa2dlwsaD7mZZYFb0hY/SrflQtl/hn3SwQpZ
MS+jPXXbgp/Np7pfNJFR7UCvJAiEUXWa95Haue4z90BE6Qf9kk7pFO0J9OpYIzh6VeFwgCYIpdZ0
bdZQHstaewR525Rc4y3LLnh8FqS+jque2sAdZ1u7dS4S82ZbiQuxSeAq3A/Nu+PNuHI7nZF6Qu1t
XzK4VYueJJ9U1BIlvhg+uyuqGI3tOihZV8Sd4OThB/u1GdJIuAUZ9D2Cxer/phnPtH/WLy71s9vk
oGUGaDbfomA3Zeif7PWFrchdj8X6nozL+wW6/LrsbtaXzhrKevxEdGMm8QoA78npTMPsUBbY1SH/
9Np+uvaXkGazgYfhQheBZcFBpQNxtv9A25d9oM+BJSCjS6eStMkqXAy5SdNAI5+6yO4Ugcxsc4xP
ypYCB7hNg1l/nrN1dm8WtA5i8LKbu2hd5xEsCRhWa2aRjGDEsW8Ov6fbSG8ni0PgtuJRMCRT+Yur
m23hoOfS7dv5QfKanuSF5r7GvxdU7Ca7P8ZCDQYG4GrSujJ0ZAQotx/qED9vZ2LYFeeWLQBxnxtE
WxcicrPGP5YULpRy5blw6N7NUo+nesyOHWESr66m+2QfcBcDaUpVoQ01N6VGKZz0GV8i528XVSpj
FF6B0Sl6Ph5PvlSmIiE2UhldUeRNlhs/KrgwftNwujYSpMNzTvS6XhAG10CePzahvyLIFzi7VQ2V
I8R3TzZtICrYpDHfuXjATkYHzZTmeNMAZV1lUvT+91V5+DmbJL7UcCH1jtM8Ttk2MG/37CyzqMxf
UbxImT25MNhdQqreueV7mWomovwn043sT8s/6JGWXCEgorDG4jMRu/U9rVdgYFQf/Yjv+R8ArC3R
vRGPKTyqKQNVh0/GKjdd465kMqj9Cw3FnDZGyp1wJWotVi/n3PhdFLiWJHs6FaCKtyGfSMqIcylb
4PXm9hfLIvjltUWGRt552zVSUKV8JzbyeGVaNHo45bs2hCiqdoNCG7nHh1bgQuCVpUgGHQKU8O7E
shdDVSrTxUK2QjHWe+OClXw0lYX894I4Z0nMzP2m7Z3uV9Ffpoqd5Fexoo7sy+dgnGxhKo8lbJie
Wte3e8f6MJTN7zpmlq0mBGiMf1E6fBuWWa8LQjexxvTF7aWR7Do1CzfnhsaZGSO09LhsB7pUoK+d
1aLZiGLMReXqKgb4lK5n534IljsV4aE2dIfU9EDro06BWibmZ6Pa6Jat18aulyxIXG8pDS0Ax4jb
kax+woFAP2ahXJHN+JFAKTPncZ4jgfQ6+2CleMauIzW5nI82yZYoH4prpqlfC+yiadtiSqewij0m
OeFFRPzljN1h4qjzjdhVHm7pyV0rf36C3/Tt6X/8Vaj7wmxupMWyUCA8q2PrNI1khLrsaDf1ZR/e
Epcfr5jOfktLI4Xp6S/lKTO32pABixBQsyiV2UGKfJGQTIJohqZ/6uGoEShQZ3yOj2LO3bZwQ0HU
5kEMSKObfEtYxqYqCdFeiq61FCWbvbTaw4yMr4HQNKzbiyHrFM64KLtcwsY86TSwlDsIs4WAYo+i
vLCJ0R9UEn8XDKNxxSs0QqhAs3LCaWSUXebQ/CPOG2O0Jb807AlB76jNZg8hUrGowiWUL/xiECI0
vfr4+SsJaQzkdWo2SgZaDoswS+g4sJ2XjCT2KGOIto+HUtovdLE+WafhXuafvFQ/qkTOYXch6r2p
pofWBphVyxveIrw4ER1GxJ7wIOzIPzLCCc3iN5EynbMrntSXwwu1InjLIeBPM4h0Qfih31r8gsx/
ARFdIDqsxJOvTLOYD6N3IivLhJ/FNtpWCoTTJZjF4MhVNSqh82Cx4l0Toia9ecNFNIkMN2a/J4YM
3ynYlJM03j3hSm4lrDhmDe8n/Lu3f31OlO7axgc+ReVK0fqYcP1cYaMkKDWgLrVv6v5GlHF977K8
ffMEk/9d7FI9WP/LmPgRp4HYKxyKn+TmSkBj25V52avcz05ZovOrhSxGIYvUbpSC/x4xHrbE7ir4
bgzSUM/blQNsawU0cT/nn4cQ34PfvtldFHsIpCYsqHLJoGLYwTBdApSUW2pR77yI1C80fEoFcfof
pu5IbThxCZy4Ha/3XXk1DGiurc12wJ17q5YH1hr0BNBQFFgWYS/xrqKl1mG+NwQce7msVHV4IaOE
WDGRDs5hrLUBECKRlROOPcSOa4Id3jijUtcxTkDcUmX0bimBrY2LTicyl9/vzbUXrIAgJoL0/DS7
qGVXl4jPmX4b7CWyHJ/ZS4eXz3UFwF4lR6mWjmczShdcFkbgdulT8Q6mnjXK7ZtKwZbhjRKbPL2n
eJ2h/gV9oTrEyIHTyh1v3XIIovoREtHMCwpUgFpiFhb/YCuvfcg/vReuICmGEek1D49X14TS7bkx
GL4A0QnNp3vFsOQvrjbAlX6D0IetBMRXH6DqBpk2ScmoWgkWAEyP54RGxMbLyqAWMnri/XdziXYT
x67Sz7XiF9YvJEUiMrUdAhc6Q4MF7r+6tlxqFc7V/yERrlMlulAhCz0UkEKRVCmrsHXypf2kM8F5
QFK3czstZ/GLjB6IuRtJwDP+9mDjYQXPYaBbDRlO9C7bPG1RZlezQBIHxXFelvdTnXS0CJ/Fx4w3
PKKGE10DcpUW0t46QUZzsecoLe6k4vt5c5e6XhPz/1433ZkF5KpqvWbX/xASO4HeckLQ4lwV1CtI
APcus6RWxI46ctRN5VorH1nUNdFJxwqjl3iyF79SxyqTTTMtdRSraiIw1SE1Zqf4XS6JSTnp+hFf
N9MhnLBuRxiHE7PS7KsJZKlYYqmhYVe2Ve59wrGlALwlGR5ic+8ijit3pjmPiSUlZZ5qRBMrwZ6i
705rkZnbmDrO72WVPTaBc0MJTRvTKAoXqtfmnMVMrkawJg4/RmVmj647pZqKs8V/gk3hTJvcI76I
gE2rw6zUo0Yyr/EsBF0vxzLr7+zDwlZwqZK971ZddVprg2o0GI5zb4PEX6KzMoqMCM4B7U3UJ2qS
EAOi1GckJaNtzyaGtBDqc8Q8TUQ2F2BIF5NKUlARXyigVXzDyf1jUSRejzVYFNKCL56Id77Y8sTD
RxVTMunSGd5+0S5j5mifIBT9C6bHsr2r4foQ3xyhxOCLScwehvDCBSnUHMt+euGsi7KLaGUCtJrg
aiM2AJrpI14PtOu7JtJUm/c1Tuf8/VOxJYlSpNFE3YXaCHALbzCM8gGegEFdimVZI265ZbIldmCs
jFP/D9C1EZMDKvVKHcZ2xiMB1LDBM40gFLdGxmwg3kRjeEDNyQQUUCuz3dUX/Jy7mJ46thBzaHlT
hvKM5DScgN90iXI783f809WRpfMfuV33gsNiTa6kgui/wzwCerCg8TEqEp5F6ekTRIBLaR4ZWrKf
7fGUBQjyogcj0BVcZN/TdcGFXDiqe9JNc0nMGlWZdnxAth3oBfc4OpErHpqf6VXUKw4mO5ojga2S
mBjAqEFZMziyoJeFKZMnzZNJjNAqW93efcQJckAJsy7QZ8qQJHq0/FuPmAMPByILYnuTiXF+eg7J
l+w09juxCUA+ShR8CfzoogsIWtzrm6ZOYNUOSowQKvw9W0im5RyjTfFMBMIUCIpOpB3GJ8VbCXPB
RgMexAECQHm8B0o1LdatLoFxSaLkib0SFcGptOK2JmBEqPYa4NRaAPxSsFEv7iZZGRSLSSIVgyCG
HYlm2oysBGfx51WwVTJH/5kcydgNl41y0UFiphdAl+FJP4H2wW4V5qLbosIr6RkZ8+ea0OccfJ9K
YHUGqySDAzzGTO4RcwV6/p8sYFZMizDoQIBNnKDK63CDwfZZQwa6vCJ/Cp2T+KPG9gpYaj4gIS+2
66tqHvHSoc7b0+VNrxQ57+Zb/HxSQ6sOlCytOIn0z65PuezShQd1X9J1Dqr7Np0DHMWKoSZlr1EX
622C230OpqhS5z8UCg3fIkAyiv4akYSMSgxyg2LpgJSXM9rS8p2oM/YLP3Gvw9Jr1iE7q48H/Q7U
icvYyZqNLPmNYNU7XMg5xgiodhvnae65r/WMdVdDqXynvVbaG4817nxRTbVky+hzVG42VD+scwXE
GodZeobYKCUQsA8ezc8hHFGm/yCZ5x6D5Ighakf0dPcU6Y2/Q3Dh0sgyZTqhpokTp75/x5zvEkxl
nxZgQKGYWt+HCjFys1QOVmg/wksU75Mb5P1XGNNcP9ByPfqbCX9NNUhmLU7QAidG9rP/ShJW+P3n
gRRzhZd94bJvS/tUiyuF8sIlxj8lB4EE/nrtUGqnLCZWTzjfEUWI9/v39Daj1b+g2vhZKlikuznY
LhbyYTu7v7/lVv956q3Av95KsEFp7jpBXWlbo0iGUfhC5c17RWUFh3dbyF5B4KiPbJD0/acQ1u1Z
Nzs6DprW7ehjFPnxlXOG4L4ZPL8xjwfg+UcNQc+YxPRpyCjxEXWeKY1X8/lE4djf6yvqAJLr3knI
7OUq3q5bKeziOontTmS3Xeh6nHE/TO9B8wHaT1CAOATcS3CmTtla9itK104RKRClWjR0yyVRR1CH
9FNgFWNf11XzkB3KUH1NvGE2IFhNo15wbzO+VseT+FzTFN/+2Jpl8+sSj6QS0x6eRBbaMfFCzFd6
NBdJGMvX3AOjpVaU8GH5T9RexWKdGUB5sGLeM3En+hb08yg/+4QZLqIjUrVMD4mo0Ap+5bSaDEME
9DRGem7Ujqq6jERv7R6lh0lPYeabuVneZfo99GuuwqgrloH0aJvYrt8nS0XAqA06zbJEm0hXob/5
7VAbjTadNlXEtZiNFDeTqXJ8WaCWH+nak3XO4QfWBMR3K5oMyzbyQV83rgvXqpE5HIALWKip33w6
PtYUDvRBJESCpHwNznaMSjrNoA/4VXM8ej+fMUibn3QgNbd3RIzD8fMKryNhDA4SJqZEaQ2dFPTw
CNAL4PbBL7suPJpso8vh4AzyqfZG4hAnuKJVg82qJjxDZorbOrXCW8/5aezumo5wzvoAsvM8FQ1a
cDSN+MdDhd7//jc7lrYotUo463pfq3OkGtqkMVV0uB9SeBnZ+oLD5bPYPZUVZZYdYp3o6Hh7jyw4
gCxtuMRUm9ysZ9XEK/dJtMH2xGClA6F5gAqiTFMA0rqFWNH9yYpay/4CR5Sya/NO/sv/Etu4ddpq
LOmuor5TUFoRwefTlw7zWoQZ2jSqgDELWA+oxWF2BGoZ8DcOOqKPDtl0NVlW1gZTlOQFIF/IDLM/
vswJ8JQG1lN2DCa7QJtRTzdFDxVOmHiGLnykzE/6nwG7G94eQl1ceAuNCqL+vcYKp2t/cOdaKGPv
MiJj1J+YzPOOcvmc71ujWDmSsoyaLpc0R+G6GMYzgw2jHVwP+/bLh/gI1RiKpxfO6wlimuSNwuF6
dBr5OYkNC+gdjITZOjxRLvgRCYxi4vkuCCFGcGHKwrkU/gtzO/QJLWXCYPn535if3U4qXxAQY/xt
PyarZ/KRz+kXcF9eJBFo/3PWF8KS/mMJ+xP4//Yz2Up8+gIuHQCTRClHuz1VjOvr2JhzdWaEHEN1
2YT/us/5I1zfqd1k8dTxgh0PQ8D3jLKpXU22Bykx3rWy1F55uApDtlYaeSjDvO5U/xu7MH4bfssl
g5wXAV6nIeFD161zV9mpape7bBSxon9myHBPThjJsXDqibfyzmytzPcrdsxiHFxordwxXbvEnwiR
3mkrWO944New6+2w5Zswjqr5C11sASXoFVSl9ZkSgNqri3os4nvkLvLgdDx0W8LTlG3beScyhBNA
GRDBPG/rt5e7BMdKtn4fULgAceQ1TRK42J4k4YJFTAQO/gMclz4oSKR8XbD9hfSf0BpplMiWNega
a9XSO2duc43VFxBkYGSqAlDsr5lJvoSa3ixQtL2H5aDREQtmv6O4yZRAo3xc9rTL60OcwJbP84v2
6VQx9Bm0h04yshFLKG8w8dr0fmoNyAMabyMXiIueD9FY36DUYGbr18/9ZaCTyx/HVmPKJOuct2C1
3FHj4XpSodRN3Ijmqswr8/gwoGfrkwWAf+Au1s48RI2gygM+FFdLrfX/CBLUFc9u/7WNye1w7Qk8
htwlEQ7kaNrVOIC/3feUzJybihSLEizF0lflkhfS0I2KAARUTBHw7pcntVIMNuqP8PxqWOrZ9THo
DUD0revEZghCfl9sdi8NaozJ8Oe234RMG2b5UQl5t9M3DIFgGjDTwbvJhFOWtFywFglq0kG3OoUu
JdTpSph+uNlkwTZODvKoL0Mw1GMD4o6kPRwkTew/q+BFG3mMtq0hPT1P4zvzROOrM6XcDRN2czRF
o+3xhHgxiY+a3gMgXR9FqEOj2u0+I1nxCCgDSkkKbqUeXys/3VR/mb1ME2jSBC+4gr3Sa/XvTk2H
sbaERuGQgpnwFS3VYx2wn4daOJ4JEhX+/VPL7v4824IrB9Uk3FhB9EnwDDBbobD5OynsPMTNDeeD
CbyinJveNwEMMpIKZnXeARcBZ7RrBy5lWS7G0mQoYLsm/YjsISJnNsytdslkm9X+rr9x+z5wkLaW
R4kD9zh3vAYKTj27Wv+JUVaFQYIaipdki7kiFU4uh94H/MF9w1qt9rOorm2XqRET4KpRKL9bLp6y
3m1mg1qPLWGjO9HjpN9U7dpklT/oVuif0mQerEPEjm9yr3gwk25bwWe6om/0RqmU9grcNo1rHs0K
zKkepEQaBr7Xl7WF9hLBt0/linaAxV9rUJvGPOJHG1BGCE231Cz/788gEvCORVwfmy0Q/xovagM5
G+9JAbGByDmLWIvnlNlkjuG0hD2V4UNBeDsqSfYIdocscUUBbtrc7igV137dwLpwHwGDrn3nPC8o
QmNunk9yPavoALPtshqCEF36OqLsuBLHVXwjjIvGo+Tmt2cPdjkF3k5nU8plMFYQQ2yYOCDB0iqC
THCn7ZeGe9t4DRvO4mL0AAZ4FJadaj3vzqXXsQsAEhn6xHWTdraFqZeqfaejTarXFMuRyGonJBfT
vuw+LNtOqnrHj05e9HyZjZlBYwtj58vsojtAfaDOyXjSy+rg11I9+Cz+5aYBIN+ciYdIlfe7NxfH
uEtJfGlx7be7Uy8WPp8SkkvNq816w/H+p0bKYDqdhPERFP/OPp6hvew1Biq1njgcvBGpsh2tsDSP
fiHjLlROTfYsZV+IZPm5nK5J8Kq30F7LBf+B8Sm2ZW9oLU/XQ6FE+OArncZyAUs7r2xFzKb24Wc6
qxjVeh16pmh2bCCxht+25VfOPgTd3DIIYgUpz4hyvNNFz7CieDGW3ePDLWD2AZjyo2z+IWz7naE6
rWMAet/rs616Gfvu5HPZW4mqCkMAyBPHtJWZz8s8tQAni+x6FbIfz7YgzMxn5zJMUM0L2up4r22N
0vkC3O52+Z+yapr4E6jfOYdS4z9D7PREqI/yHAuYlTHvg/ahCTgzfCWvgji9emEMNN5pc0+J5D0y
iLhWn5/QxyLTVBw6MOAyZ7nwnrO8hBxcTE5GW8RFe+yPt3wn8NDw6qJzxLMHQKZyOqDD4RYM5GKL
RRYB9QXdXozg4j97ZWpxVUAhlsqRNayCGONkNWZfm5chVa9BU2LaMw/UbYyfuxyBxuHjlAkfiJ2V
EguU1RY+ev0g1jiqSkEGc7rJoO6Ma/yDyWbmBFZeY1CTgwpjJ97E5peK+QfW+ZX1XrFoRPS90zCa
dtaG0ewC8dZJJOgrmjBI8xal7ioLBqO4WESG89Zp4+mhf4rOteeCJX06CnuJx1JBg9fJHGkjWBme
Tov5QQt6aQJZoJ7nf1I8T31ceJU25kiTkgnFU79VufAdmJ4Kbsr8iLXGdDy7xAl3pQjcRNbQ3cfh
nBuiWE1Yh3X/Tjp1oOJ7iklChQ7L6K7pfW61axzmkE/1jXnRMkDAglN68JMlg7lCMF4JozU8YHwY
CvCaTX042ljPouomhS3kDcsSigWyUx33CZdt383pGGUb4QR6KUJYckNTT12vx53ZiZxS0z2Mz7EJ
Q/rxtEOkzAEqGB5P2YLGqv6+EHqN5EIesQz1WaN873GAMQoVqAJTBPTA1fk+/ZkqY2E15Jabth/a
YhJ0e8tCNHprbz/pByfcb2BnLi/Y1vHXJBhjmaJxEE7kINg3KKr2PEHauTUdTNqJGvqLzECkkbVA
wu2rsAsknX7eq2xQtqkr0mRJsb8sOL1p7fggO4lHB+EtXjnJSE8lzZOwHcDTVMllf1iGOCjB2K02
L6oHATl2K5aRZgTLzkSRZgZH3BrcafqrS2nXN079VTcyL2VxJIzrimAAZoJSb5BHTxjnPaL4ze9b
kww+oHivaOxhiy3CIFLrV+pMjzkqpHfuqyN1/oGMqM37IF40pngwWT7WgHG4ejO4qVWTavKpOlIw
8kKU51oCmxFMr0b5qbTTIJIhL4aqvj7/7e4nmxTh0I9XmczPk1w42xarUfyjx0VwoeiqKox1osCU
MZI/+wrC64NLvuD1nr+A54sJdiOXH9nymXV2LBZZgZeaPth4zZ6bijOPJeOHnPEL2PGxa3fHEkZb
FQzD/53sN2UFeCY1dv7aW3RQqTQr0ug98NYC7HnYTlqh1mQFh6nKZfBgtQHQOUq8V1hwR7wEyKBJ
ybnY6uN1yLf0X8mGo4Q9jWoM5AOEKn0FSKwID3ijmjAtVrLbpoZgreVo2MjF5YllTO3+vOdR74i8
3EhZc1aAlMMjGJjIsrw3YtKv4hbKQ5XydS9a0fycT6kc3I7Sx+gZGZ4uPBu21izxvl/ubHXhNG0q
deyJpHR+V1MVV/LWISDqLm40Xa5voJi2pzbLX+5+rEpKX1Uj2P5zADVL+QVlWI2wLYwS9rAR/5VJ
MUNF1QLjh6J7XrHTzNQsZ2gGSzO4EQSaUFiMn8eqzUcTutiZrdNLuNZRE6/JcJLFYdEYXIvsiYWF
12+nWhoAk9dM+0q3t3Z2DsYSBxY4F+d5fugH+8iVs+wEfkAigk0cMABNnQtOxjqWO+/P6bI4YBRF
DgsUhvOQqQGiPdvMsjQjnKoC/TG4e0h7rxjKHXSW5uNJbCU/J1OTpprX5MI2NFksUXcT19AR83kN
7i1IROL5WZRdHSAJmo+WZdhKKL5GVPU53ujbzyyLXyBd1NMaE8jFNNmjW4zMR587VFw7gbA8hTVI
MVtMs6RclQW7d1otX8I88ki6BJImUj8jBfSRRFrqmo3wDaz7peF4AYzwH3Yiab4yG6rVTvPsZVEn
p8K2Cyb+9KRHTXgjGnletd85YpKxnh335A2b0DuaZ/3qVCP4BgZJnuPcUS7ZIxpz3ErRumuecv0f
wlyTAeZysX/PXmPiS6BvKyX0dDKpPBBk1y1SU/9yP+2+eaZ1Hg8u69vTIq4nav/Ms22rB/vRm2ql
ZQh6jebD3weZ9y27PdmsZELQP1bZb2GKxfohaQI2Ybh+d5hbPukCjb2mhNF8E7OFUbhEJZdWgTqX
dCN4VPUJarXQDEW8Uc6cSvRPVETmfxWTzXel6N9RryXuO5vzo8sDTncyLeBmhvA4NnY04ALTuiJ6
VaQEzYKpSufbU45tt/j46gm/rRzD3zn+R8l+0+1VosAElC4ihNE24hR2+EWH/Ga1qL4VRzozTGTm
BMLi0Sjjzh5BRCbRm9eNhTt7wPmX+MI9YpsjYhe9BjFbllVPIS4pekpvbfxCNGYKFmhBgOf4N8yG
iVqERxL+MHOxfYXb9mY29wlErIe37iyvUNmXPgQZv2bbVQ8uwlexQMzee8xScXKFkklsB+7l54P4
zoexsjr6n+PwCUDx6SkOcp+EFNVkRy9rEcyAl6oYK5DsMyn1QqXNWacwaHfibaiHVxKpHopoZG3f
8Z4EL2xyA34kPTpOESKsARIZIb1maEtOIUjBRl0SfWn0prUuL/Fv+8zD5F5MbMuYp6pDG2FeY1D9
sDXqq6Des5b5DF2HCp3ZyAb4gw9W+StV/rRwKmWuML/3QwXKu3D7QngInCh7hE0WoK++8WizcjyR
38+uKtce9lKTpRDbA8ZonPOUTzqUWrdpoOT9mVlioV2uy/eVNUECketykmZDoxUX8OGGYGooBJEA
08mP/ltMHz7fOfJLnP6Gx7DkBH4BzzWU5U8Q2Rc3n3mlWTTpogbEzk9pRrKojPfkbdUUmqux0ms+
sgTpa6ASKvMlcK1XZIaDAQL4s0o7jlk5sB2gU5hZ15CWzUKFkiK45L8W3EEV7p6dIz3Xr8TPFZDi
pBp2jA/dvpJkEDRJ7U6Mkeb6chda1II7cZqlWl6pTFEIep48Q5wF9FAtmlgX49XjQQZIZIfxJLf7
ANdfAp0pIQjoIzfOtYX1iGZjg9+HO6z5Ze+ZMyVMMYFxe+QmdvhraObB8dkp5eIEVFeZnUte096S
0fFhWD03it5qeFZAlk/XbROI3+nqlfli7W2mBcirhBvdbtfBNWAaAMbuwaRCVVgC6VYL66lNRTH8
meLMJmua8op7WslUbUGMo6OFeStJu0Ezh31qAZelCoqIc4a5L3kJlw/e3Ws3GOXLh351NlxkUo5F
R2CorPQJZ0ytnjpMFdOFpyqcWoKLQT1APx8ggDO6Ix4QE67440SDHYsZq5VPTnmwJYUu4n3q23on
JNtZa+nxYEm4m3RPaKDTe9au0UO0X2wMzbuDJxb3++Xt+7RsqPE99wPD61aijnz8K5oncLK0RoVq
vosnr5CM2fFJ431BsMhZALmGilZeFrCy/47cfXawFNstNsusAWI67rG0GgHRkBF3wIyEGotgtpQJ
SgXeCeiwndzs8yz1igWWGmKnMM0ieNAn9HUNdv/vyocaV19vyGO/mHwJAk5QrTdiK9ilk1FTVt65
obJcSEWT9SrkW8MmDG/iIzdqsqX94fcJRL6/AM8+MPCRFr1TY7/KDwgfFS+3vf2tYMb4o+C6j9xA
X9GTMCfBSsxo1KMuPBhDqgkkMbIdxRUUtJe6zKnPvI+uTKulEF67ENGI3F2w4zB0qREcWd8clWfS
QBbWaLaNZ/+DYwe1waZhG7z1+rrCZaC45MPDFZA7GDETC+0MekuB5AisGsHPCcSB7mOg1VS7Ghnz
qkjBtCHzt6PJT3D3EnZi4IYQyS3OC6jwDCsWmVz9fah/ulsstTzGhQM4zUpfq3spqtlLftByCoZ3
R0/dBdHPLu3r1AAJ+6VGsocIEiW6hJurY1Bu2kMRCtwq/v8MaK5bX2IqgRoDGZ+S4TJnbiUJ1Sxj
qkXxF2GZAvesoaFPQnsXLgx4IIriuJBUJpPsSFHuH8DYGDq0cUIC8QytjmPVqHFykMmQhvLfvQdJ
3Pgl71jBIR6+A+pAUxqokBYQ/9YACiiIOVzyycjjmpZzUH3k5qFiJs67p8F2M/ybmrT4ccIur9yv
4wra1B6MlCpmtM+VB3ZU/0T17rA5FmlwJMFYUf0STGmrRH4QLyEct17IBQmeLmEAZhVMPEwkCDjc
lHJbI2GnXyR/EpJeUW/sQJMqy+VTPjMF/JJOK9oGEXf1vqgaFIfvjxdebYcX5DuQFsk9eicMs7AU
vO38HGG2SHtn9Q4pjG+/Q86ZdDd2bZ5xvhybwuPajiZ9XfnyQW8RhYJe7XtwZqNlK0qfwAxERemR
rbId0nxxqclmnPEIOU+DvnEhOTCNDnlac6zQO0kBMeSeIaiWgyxXADkm+QJnhwJ/hDHUVZpOZn3w
N9zzpmwik12rqA9iweYRxqTFLuvTfJr4fzzYC2kBf4Cl7cPZN0AxyZDmTfwdd9Mjm3LxA/Fa+9fJ
f7RkG3oHf5pOXaPwj+OzYtNITJXpNFT2qC2mzNlyj1ALKKKH1IpIWDkKocAvI71XFz4ZHnnSZyOV
qaNTfRl6lPViFAF9eVy/xvCrWM0v01DhFO/m08Se1+AvvNVJAbPMivLpK6A/EVWK7qfNX/WQL1z6
QFcL6DRy1V52rFXU4uDSrqsX4V/afn8LAyoItpJgstAkUlmpXGfPH83XD1zKovXAIo/m4+ag5YBg
jbUi0szPXnZkHXO17AR6r2Dw+/aPYDHYPoljodpCJC+hzNHjRQOrF9YV9H9ETcjLQF8GJWmBjJee
zJsC17l+oZZyxUMjRNHHc+iokQwYiLzyybds/1xQ14izAs5Jwp3AW9vsYSYq7OeDgKwtRPwFVNgr
1W05gsdI4+apl0gg4++P7qKktKP1oZPchOQWkHUnE3UPqovxEoM4G2SHU9451rkPv3XImUQ5JV5p
E9KN9gwoIDAuANrCQ+/kqqJEtXOKQCBSaB0yorOCfTpT3MfBZkxqZKayJrGqhTJblnNDaZcW22Do
Coek/hp9dCKy4oPbQnsjsV0lz4lTruV2ybnln2LUJCPwXPSatC29HQgjNkl2frYOWUDEBlVfSc0O
GJRSUqjPH0g4PgTruqMDmrN6NI8DGo0xlOqKTUuR8fRQhvAmR7uKMh97HtmAGTXuEpGVBkS8kcad
5FGv+p3uoYDCXc/HB5yAHYr7BT/4FYb8Uo5pwznLcEYHYLX9u2zfD2dKgOj/huqJ2jrnYBOjzaB7
z6TiqmvH5JQRd6vqDnjIeu6BW5LYj/XGSzajqGs010bl4N/2IAs6sB3tYyySaQvhJtpEQOq/E3go
GtoVzjaucEuNNNDHqhQxieM1KIb+WsroF8k/RQETAJu6ot+57GaGuVoLv0ypKZGVScfAcHz4dgVM
uLrEwwSDQwwQEMrlRQn/GdZSVUSVYInURqC6qtFOZjq5ouZLCXh3KSqX5NUpqRcSPb4GgmTeCXH0
CySCcNGyd/QLtksTV8aqVtwOp5gmFo/Up/kZZ8LKnYA9ttpGRZUL3Gtu0HMohWrqqsaAdL8r2GN7
KjwL5rj67fOHXvZC3POy2SrEvE5kLrL1ph0bsKU/lKa2pR+XfeETANNxawJvHotYUTMZxIqUe1jQ
R3RUi5d3mLzTj3Kl9kMbItxU95g9wA9z2qIIjxRJUYEebMCI3SZ2Dp9N/Wax2fDzAoMJRGXdFqsz
BtfxZ2RTu4a0CsfTykUnMykzMJum6x0HQ2lz43+2krDWk9ivb9WO9/vXjRBg7MLNsj5PxUqOInhb
zDusNOfo4aB3PiEZEYZ0XX98D5GyCrWuaV8s/8yiTv11D4VhF3YiIFa5UBJiZP6EkbmRPAxMqBuf
NwFBLR/IdDagnwCnpMEnwCywLljm0NBFDNsbJqWR0jn6c07kNk3J+ccVGOLJxVx6ZAn7gjC30KFz
CzeLH/kRR//oHAZhyP6LiAmycoc1agfcBMpMMydeOtfzlARHekQdKZQ6lBhRUxB7f1DCbRki2Eex
Yio0eJ/Jrp0/LzqygfeTRkAlqE8Mt65KrWCMZZ+c5IZTrOgGxEoA+An3ueYk+eQ0BXA73rvddmGY
aus3yWEIVYdlnEMi5teeJqN7VKuTXM11l5gDdXr/IkeopN22eL44OEymNbfgsAySlt77RIUTvB0f
ZH4Di9Y2SHPbZ8BF3Mi+/PBqPq1bjxXOVjfKzroVStYyxKhFs3uDwRkMkaHi+AyHXOqpsCEReNnA
Dx/uv7sOFcpQUs8I1QhqXLnCL97KgD9w9E0UtKL/ETw09zYGHX7ke722qXWtClFgJgmNqXdyf5dC
GBZ3l1mEKUA0cFcZ2gYqMP51w5z1aPTcaRZnAwq6QPl63ycvFcgSoVPWSwU9QYzRk1nKmX4DOHKn
NSeb26pgBkK4kB9mnZ5q3KQE77eqLDHnnWngSEAZJ8kuNEwjs3RxThOhHfcy/2qIP9dN4qjAp3n5
rLnIKOziNQ6/US1IMks1CW1IkB6XdY5YPTrBuB7tc+51GNG0/99gjciQ+tP6sWROS7QphKJzjjs1
Aey6dI7oCZL/VwukyWndAssjLbZ/wwLa+MRkm3+1IJvwNRCeQB5WsfJrIU+vqw60I4IPyMuFBmbg
yaTUiX3DZxtAsODGUvnZq/iW/7+HA0mMIRaXH8MX+9qscUt+FiPVXXczeoX/yVMSwdjSC0KlVv/p
eR1O5oWibZXmhME0PhU4rwma2BRwr80W9gb76HzVCjuCjgUSYcEujTp8F6ZDZHAWcuDnF7XSw25u
jw92fOxWYHPkuEnb3mD8Q/yZ1jKLjYz5QHGbIG9KA3/mS43T3c0mXfeiAYB5eYE44USyZTQByaTH
Lrf/I5wixqMjZl4yKghJowIpgwZujqOpZmDvWw3Rnlf4F7iZvisaiFN7IZpZ5MRAQSX/dMkg2jJh
roRnr6yP/a4u8NSsuqonceJs1aJIrI7tFZTZeoAG9EHttfAzZDTaK+JtegHHMaYdbYdatp+FOG74
c5mJK3Ctvd4yUT/DRvhK+nChJFg6bEcV06OU0BSA5U/WtGIGhCXYkSAmga2a+TuctiLrD4U0K2sj
Wn9IaDgDmTwoxCdyg/5rs/pirsSm2WnxzzsY+SpB2xkDNRj0us8vpv529KKC/Ag+LgDcbJMc2rjq
vyZ006jG7U0ggflewc56RSFx00gohr9uIqAUPqMYFeRmI8/phMoXgCXbSsyuHdw1GMz0CiTx66fN
ugRY2tq5NZf9RSATY3eZcAe6TOY0pgW5wp7EVAn22tzOSI036JsCoueHtGi/M+PVSPOE25DDdWYy
43ei+ctWPIGu0Of244JBkWcMw2A9YCZK3FXzsW7G+fVhS2+Do0rz612d6lFa+sV4M5MAqR/GRNd8
BTu2BPrpSrd8O2SAV9va3rNZAkVTuhWw9RFnNi1jksvPVX/0zB9XTFGDarAp0lBrj8mlEs5vXDBM
dwj2TsPLXRIkPpU5fkkcGW49fw5k4D3ZUWQEY7rG1hYpejjFtvp0dg7GQYMB0tFCw4MrGaqw8FEq
JijeIsgeKFxpWwu+fXHhpfj0CAIBkGrITTLZfpopc6QmiJUiTVyGu3VU7Zqb/cohd3PpwP35uGK4
BBVtx+1GG2UKJ3FQe3X2MDkXDNqrdCdJMuGtTr7nfFE60AJSNFiEHKUUzpSMjzVvOF0IkGINqmAL
yC3BTzu5wDExj0zCG/KNHN0VMX6Y7kKoqEdvN2ttwWDYYQ2EOJ9I4vpFjDvs8UZ+PSieaKCJ83MC
BHvcGPC348Sscl6gXUxX55299wB4l3WGPLVJ7jWB12/gC8R9gdlYXEcHxeCO9yBsBYwaf9IqYX/C
YI/cdCXBqRlfKHZJVFv0TWz0sdXOUp4Xb5ia+4p8myabUr1qXpr58uh0xSS2QcDvL4R1tHyNy/u0
sEiviXkirrnbl4qr2ex1Rt2vPNgiDsGmGc3GlSxFl7e1I7SY+ing/tytcEfgYB+OZohS2yXLR57c
mtsyA12tb7hnTBLjqBzZsO2MzlH9Xn8v/PfxVMTNDQYQbDRIfk1KnqiQM4FNKgSslofjtIY3fJp/
xPQDkN738V1dc95adZMUo4PvJMGWQxMuDXWT/t5CewP6RYn8j9G4TP5EBwAS1D56ue7f0OVsKAGl
njD6OS27UkkgHqQG0C1SSORu5aMYsoOIO8OWmshxhkf7HR0gusfx/pUNwII1wxNNn97GLQNjCrFB
zB/zfZ8WexiJcAgBQdGQRHileSLIBA1/iLTv84D7pGloQGkXaLev2T8bXgj3VCklyeR///P3DCxX
mjeWIGCMdy4++kB+M+MhJqIypjEbZW409Iv0hCaiVK0UDROFkV0QGzSNfE6fmcQ2M04p5H91B6FD
nAIJGcModl/uF58maICdW2npiTyOMqsc6riX0SfapAUqKfD0Jr9ootI75gMZba8kJM0/pdMdM2A2
xUUTT2c0mLLMDip8MerAW2KNIaXqCHMhu63DyrZ+IlQdf+Gp3y7E1Ejwvo2G+i2FvdsK4QJNhdUe
bMKBYv60dsOAmVv0QNAk/sTvZQQgUhmqgZ6mi4+gMDGEgshVsip6fWoXJjlIiNaPDHlZUZNbDbEf
OTaFiFJkHYeRmxPYUAoEa3BbhSmkYGCXQHRmBZ9uu/CRGo8EtYHtxLt9heR5ND4NNKYE89iqTaeS
HLU8brD6jXoRwadkYydMyazuqOuLhp/qdQ6Xfedga45NMdiKD+nxFgRb/scZOXmuYkJQUmOoC1pd
YXufUGscnogsH4GKy7tsd1gH7A8IQQKWGF/9YL9gR7J8iFOyrbS85XtFaRxc2mcaCkbDUV8Au/Jv
q0qsgq7F7YS5dvypyHqA50OVoVh7AVR+zFzpnW2lg9NNxmcSkC4CtJ0kbzHSy6y+mKI7L/6FW8PQ
Jk1N0Ln4Fh/i/0cYbsFsr2Z8lhxwYCYMv/sIdN6LxZXWSQbZrYZPD4xfZOQDdsarjhGnrXsQiAZI
WZY3gNwQVJ1aWZbchT8Cmy1EPcXzul7J5KA/G/1yGn7beYqKMt/0i0kmCBSI+L91MDuIO0JZ/ahE
ZrLAlcb8GxDM8FEFPQeUi4uaXpvvk1t8ZoIdZXC35tSQiSPQcP++mfX3xLK7neXFyVX82QQ9o/10
mOwf9rrfqjj2IYCRcDTOI6pjqeUxUXOLdESCH5kgwdrn3T1YAAkl9Nw1Q5c2zvZdqR9N3W24nYaY
2f4ll2WyZTWIQoDyjja0hqc2nm1B0vnh37yZSFkgvafCu/eTRU4Kylve3VvxqZ3Ff77G8rXhAArI
bQzB7kiuNmtEUKjGiP7eRhsTMMEf0d/2GlfHcDztqvzyK6U6cfL9IIHVFsjEvmD+W4TUKrFFhKui
Hrxm5zBVXr/H9/W3T6X67Fy2KyzZWKYtBzBEy3Mt5F8RyFjYxfCpP199CGXxT936phF2cD1pDZzb
P3buBFuyobSpMgbcFV6koC3kLSJaIzKZHzNg2+sZK4sbytbVjMuxDbR8vYb5mCBj/tdWOjLBPgrr
c6cC+wPUWp5GUJtR4QeE49Hg3J5HJyvCZMJdZsDhIlGmA2Zt+Cy8tToZHTVmvHiUGkAD0zZT8XDm
cJrBwsS1/+gweskmaCWINefqAaZQ31wAmG84uquHu/hr+pI8KvGWAQ4ZejpoNFb0ulsud0HFCHfO
Sp83GRDWxb5hKR+yQXjASAtqZRqA5HJUBUWY2d1UCjxsLoQEd3RtUHFXaxrgLEFUuwhVA5g+Yxmb
Ef1wVRk3pSRbKzQNV5gqSkrFuowzK2AVrMaT+u+3NnoztutRefZRZfwvWLVe5yVtnpSRQ4RIRUeL
g3gggC/mBPalYnM760f+sJVvt1eMklrX6RxAIunVFjyiegjTrcbrXwnhZoV2UBsWJKBg4p6VFfpg
C0OkTFUZ2TAp5t7epyH74qevExYnbS25OQ292jlgL/BYwXOrUEWnPAl+AcVNo8XchGyJuLYIihXi
QQQmTW8pRmAOqObFt8OM1p36PeoQISIPXn0mKQRt8Ihy78u5+T05F/LdVYCO97vfIds4n67N7toU
A/i/G2uAYRWvBkXhc+teV9PL0u51oeqijqqq8CYnv5jVTbRob0d6/lXPKtKZm3rVOfsmyGC5Uej0
4450aGgwqA2LJ+h9OqWBVSsaquht1+Xsbmv4Q1mINbTaAPoxhkOseKxeTbME+RBVJTOtVgcBixDe
GTIqMs1OtMtwTL/pzrs1ow/exBsNpN2OcuItGh1/4LRAsTY3wHxUknOPC6NAH5wkZ3zEFH1vop/I
BBAY/PawKizhYgOXxZ73zx7P/IToIli/yBbidiA/pCM87pMEesNEia7LMVo08TIh24wybZzZuKPr
RB0hRF+8EYOi3f/Ei7IvPT7Z0FciXYdn/YLQXUB83/CTpoQAJM+NNfOGBswyVQcn3Ayq9GqnnMoX
L+yLbocI+NGTuop1UkRayKilHYPrk5iiiSp2J1iI2OdulVuOReT6c5XFhDYYBU1QIJK1nqU4dt+K
P+AbI50ljM1QlfDtjrMzeoz2rCo4yc922M5sKgjlABKSoeZo66YqQEbx7IqNIqKA/2bh4tAhHDgq
FVLRrLPN/XA6rpsdwCowCXcOBn31OZ73LIisto98iSxAqL4oagEyRersyMaP2NUmmCNDoD0dT4oA
+PGvz/6Ttll3pNWUGWsMW0oT7kFxReOE2gGnUbKjQ6DpgflsBh39Pu1ykpNaYoFWgw6arge5tMdp
Jhe8DRNB4Bc1im1WlfFpQL9v7xXjtMcCuG4llUs9/1UoA2Dborgn30FFhGDAfG3UwbwNIwMGf54a
mG4Zo0V86M7A/3LJ1B/w5WLds5umoE/s1R79a/joNL8rmHgDcdSbVy6GA6mVTNQMtaetyiZg902t
NxFIAQrzBa77Ax4y8mqomKHFQY6OEizm9pEXAK0zvuanjGBws0tJ8g7kIA7oZmp7cCkqtLMvWU4H
WnWw73pa66nr9IZahqMr35oibU5W796KxnW9+JJIH+2RcXTdaH3bTzDuz4+rMyMIVoVErga4pSz1
HbHfXahxCsZhnb8OU+U619TJSIVgRhTpySMMG9BNA8f7ttIdvSnNxs+JgLxxAsvkL0w+wDMEai7P
nGfRCeqf8MRJt5sxbiYRkzIc/CKTGvQT9ZvMWA3hgsx2PZplY/5104ZfIFugeUzUo5UdrbIm3N/t
NTd/H99PJJebcx3cY1R1LLtXvJuKw27or0OVTy4cPuBhvuCNxb+YaoYplwR9rA6fH5acL8bsHm1K
XXYE1iI7j6DcJMFfGmIl2fWnMkrSqWR8V4ACMGLgOD/iWtelkHzvwSKOIovm6jOXKzcVtWF/gCiv
r+iiJPfb5bCSolU1Z8KMhUlnoCKtzCkuiWFPpVrFoiPPPL5rC268jqyFESZfCnfbEI32Su3NLUGm
BqNXTKCe5OBsgWmflTk9WM448duJLQh2UU+6dWnt4XJLG+LVRClv4fSYfA6Y8x2A/Wdr9v4slodR
pbxWXYAwF4kiotibFKQVH67MQyGwiVZo67Mnte0atPMo+68yudQa0/rUXY4gBD4tulhskz32PQUA
uD4elTXDngdhqPhnVQsntzTqfl1gJB3krDdl4UszC8/3EM0tMqod5GWtuPbT4aUUZDjDf1even0I
hNc6xRPLilQq1da6hx4AHq4DHAcaAY7CWS2hQzqTINuGqOPSxBqX7mfFVhxujNlrQiQfcLNcZma1
zizHKm4uZ9q8h6FcJDFDnb9UzA9du3auhh6SDXLxazZtKKMclmJ01drSSd3hEE2dqKWL/EjWeEv9
7ATOzxSBP9/RYSHhQhtrAJ9Nq3dqrk7l9Dg1ORU9WPyX61l8Kir4ZeLGjGFk36X0O7EI/k88Yawo
6TW94EFVWLGFSuDrDiW/Y16srLTGyWFKqxDQj49StyzyQb0sYKTzHFkMCqrm10yrtSal8H/l2tf1
/yudiIXs04juLqWBetnI6uToeFWuuLDVx+3wQB3lxb2WwVaqEd6cNAqN8JmVbIV63J+Qd3Dsm8Vv
YUFfgOyv5YWTiuCtRfGGdStipW+RSLQYar8ggs3x7zy4Y5/yp5e1PBMgedf1R07wO9e9zDpuUMeR
v90VR3/pByHSTCtwnQXK+Wnq68ucXhen6AqPUIN7O1lc4tgs3yMplQWjTyuau/OIdva/HGX+5fcK
exUJqpHgqxnkzIpqrK//7zOkG54AL4p0P9ZW11ZnWfw1QMlFcDUqkvzOke347ATwWBx/dnrFpYs9
SbJHNPasWgqLI0AKA8pYVwDj6NxhmIq+XCA1M/NEPbkEbjj9cMhcGF5HRcX3DbFgZJzeFtZgx1no
+H64E5+7tORnLMlA+BR7gcOIrq5n2ZiTyTXMwwlm4DzcUSPEY8weo0zWNEb6X3K9tCEjGtGWxfDn
Cdms4yjLCyHUTrfCQpFz5oDcDlJqO3t4etMLp9YubuDLXnDoA04J5wUZlNUdkVbwXbAQRjzamJdl
NbSEEs5mF6+mW3TdfG0+pa81viaS+4eTaICt2yCc0n/W71O2S/7MfQHARgFWZPRZM71PPiGggUP6
tz7HG3ADx4e7VD6P5HYiEF1BjXgzXrRuo8jrTwLDwju+B290A/DIAxJjsB8tXX6Xi3rvJnR8OP7v
zbmjF6fghEAYAwg2qK9MdIuJCP2lzGj/hmsam+6YnbmOGTruwwPv0tMet34YzX/SIdS3err/6dym
AbQMr96aS7QPEPu4IUDHu5flJW54UxQQjn2jIHeBZG4PbGaIrBIpx5LBAIoHAdLKs/0WI4G9kzDf
LD9dlXhiDHZdJ8o0BOqGrVO+rovcTg4ycM4IesddocDUNNmBTzsH6WxNUJdDLeT6J+p7h0xEz4Fq
IwDbINcxR67U0MznTBuz0Z17Be/wK/K5JWHHHOCnN5udiq4bV9Xn16+WFWO/bHsgxYW25mkFX3jX
P6G6vZkBtO4SCQrYs/7SUck8KHzVNtbQteV4ZN6XVWyj0A9U1j1tV6mzBS0Hfomf//df2MkcO/7o
YqUYIXmKowjlsWBACDHWD1cPAWH4/pY2CzPSWFB6dZw1sDPAQ8q2ZurDCjDXjeQxzJY8JnIONExH
TD0fP9Hrf2fLzSxsNMQspVoZQoIWJ3hNdxNmMbUaDP0UuAlq2FaO9t9RkhXbv/iLXDldskXlRqb5
vPwcgkD+kAQJYuIAt8MRAXwrGcAK8b8/9uv+b/xsWxWj4CR56yhMlvEmr8urCspTtpoEjYr3pYqN
k9xJIQ601tdSeQYp5IDhW5yS6TZkxL6T1OWrA4qoC/Y+wIf2/83y62i3qwz0SHng2JHyJHy17ie/
cEY6grZOXZmSUInU3ZOG3IFsm3gkWEfqxXZTiAL4klOTN3rYXsqPfxNLm5NkAkx8/6wGwlGgOAX0
Xok4E3Htnn+QiktbO0H7AHCBDjaB+EIHKnZhpEa0yxE5sGcTzWVLpheHMExnN213uukE3mxgHKel
rU9yxwi4I8U5NERYRwN9ObXH9+acg6yFpW8+Px2pfRTzux75R4FxbFBIWR5XQSTYMtKYKEhZcTUi
J4bTmiXFf8p0NUPMQRUcayJ3yILAeFBm4tNfyVKlOrDbf9FVBfJb+AftV6Efp3tV1BmF9/XwMvXr
8E7cjVZvNxKmB9lwx447y0yFVFWTf1sOt9f3FLM4nALFu0AHFh0l6lOfnGeEGLOwctuVwl5pUwe/
ktzQDjkuIlCpcVFr2Cfr+XLehV3GNG1vXsexM/3DyUGgj/DjVU5tY24htp2peWu/ikutz80s1pyT
xNaefM1kBBLjubqASvbnmbrHwK3Qnl+GVwt8ZR8ffxKpALWZxP0Yt80b4nAQy/iMYZBp4ivqkDmg
vVJ2FoRCZ8bn5kNQmcVq+xCQ44Jo3pvksZ/mCUJMD3PyxRcQFMPXVlMhZCSGQ3BsN2fFrrG3C1xp
lFb0w4KzYi1j1rha9a7nOmmnF7SOa39RrhqHPD0EjXvELWN2YKlkonWg8KSjSc+sTXSe+4ZHq8kc
mnOog4KNt67H6UXWRCODs/2OV5sjG0QbCLtXBbls+DHwBA2NgFLVm99YRj63VRRN0mmcOtFRB/YR
GL9Ep28NY5Wh2Ltzl45TFxJGQd15yHsk3/p8Cfb5cHIpMFtGXmwoSmCp0aFGJ0SPwElfbNLCf4Gm
eV3KG8aNZwn2kbbPortcQPr2Ltl1PG6y+9clKt47YjsgqD/+u+90pjKp68HjLYvEx7WD8U288sUq
PxYx0RqLLSRLt1qoIaE0UwE7Y6S7IWodLy1IkLlTYhPcNoyjCxY8j7NE6n931dhME3GbVcPW3a/+
Er9ieBoYIkCxn5RhTpFgxgulgg/eT4fGbA4ANGkJpto/INnS0kvWRYjk/KFDo1YWkxgdBIUv3XzE
c46Zr1Dxq7VHlAbQWzyAhufQKxuDRs0GPFa9XPcw0cVHhGZD5s/kP15TNqec4TBbIWmQaw7AGzqM
J9+YLI1C+9riKzUP4d0Fwy46nXdAq2UKgY8P1L66glyIuTeWbySP9JpWjHuagEhpIvHAcuXSTKxk
W6gjc4xgQrQdrry3pmE7/zNeWMxV7NPFn+L2xWLqa1uWqwS+0FYluuGsNaCteczJAtYK1UjxFsMQ
zKvSOMnrSs8RiQLZf21eVMNiLZfn0djVNms7tzvIL9Dj3MTxDSc6I0ISIR9R78Me1FLxzUfHC4yq
1EUh0O6Wi3oCgHjUhy7mip7IDNmTqRdHgZeF2OW91PEKyDjb/Vt7kOxCR+xuKHJGqG9tkkCd2HYv
YxprfTZ6A5kJbFQX5W8kqZFhCWljFqWkvBpmnP+mk0mVsLFeQWGRUQ4/E7gYj25+7azn7ctVbQH9
VCRL0ylpJ3DJcT1OYePUXm8CuizvvQxqhfd7Ja5mFZpHyAo7bN8I4jAgzPBQuJris9B/8yf9qTcY
CzHiKlESB3CdJpovdDaG86cwoeRbAhv+mAncGdYsWGB6HWqzxXXinbvUbMUHihL1l5VdwVaK/lKH
xfPM3JWnbIA1ccZjS5rWIdVj1+GhMJEY+5hVJv3rHRmnCbt2KdLFI64WyM2tLHnelz2F8Gns8nka
C13Diw8mGFWCImdCizsXS2Io5KVRH/deB1cVa/3pu8NHJ4fZis95o6BJO9HWM/ll7u4MF+mpFNnw
t1NXkxw7MVnywO8g6n+8UqMzjFtt6uhP/gubw/8cL8XNxNfP8B6yY1XzYwUkzvuHXWhx3YLic8nZ
pHpIWbLGTTFgubatwGxsvAzmWOdNS61tLmdGuO4G7EeKvMuEeZElD2/auLfD8PIfBOfuCFT5DJM9
zKgHE0bLtpuruOrlxvH+IKAilX/6oEw5S9IQVYI+G+hdNlUBqsp676zn0Ok10iwP5igNZWG0MRiS
2iKjP36tsI8BY7I6HMQMqKieaOk3iOT1M9g9IXj3ChC6yatg1fyQ3vRcX9zEQW34SYoAx5VPP/Ho
NMsonBaaigWdVegngWlprsE/VWFum+wL1kim8HJ9hyhtUtl43XQPaNmBurqtc9u9iL4YcJtS1VT/
0H04XuaZiOapHKj+l3cxHq+aaUYTA3RPiQiQdZ6GgzRXPnwsc2t7wPJn3YjigBfnJ99v5CJQfL6u
O/vIN84od1cj4b3/9GpPkcCaG7zcQVEGtv0YgNC8LwwaRB9+DvDan1tvxveSF0zG62dMnke8p3MJ
rCJl9h3Awy1sm2DuzrJ2omtPXnD77cmnZwKOzqh4E443/wYXa0BfzF1IpEJJXZfviwAFBWfgAe4r
vZpLG+6vjwqcOGf/MamLFu3N5JCXqvpZzp2JIgULiUles6oy1Bkuw4JvwXEoDBLMbpxr4oN4OURM
4PREZg4nd4Y1OmNQe2LxxInn4ffqyEABhQXDdCbNlXqyiGY4H2t3wRDELdnWzKS4JyvrprDgGCyC
jFKyX331TxOos+0k3sk4wTgwFkdb7/93q2j3Yd6C5vqvXTUqAfTclt8gLKeBULizKj7Sb5RmlHFU
4NuXWn9Y9MBf3jRC9ia+Pu0Fl6wDCmhgkxF4hCqw1chnwQSCCqp9p2+4I4F6F0QxQfbUIN9HPDRk
p5aPLq2NAbF5VxYnEdJsQf6ntap+i3BLyn9//XMat5vFxIpbuexmX7FG3nniD09aWUMvWDfs0MMD
AxJN8r8YfB+9FaQrUpOGVP3IkSS/xKMpoezZmZBk8JYfyftV94UDkjyjRGcI29uRWGHq0tNfm3YY
YEeZ2r2yU0P7822t7iX3BpDUmBNvjd11GQ04QhJ5ZLf9VIbtVPkmFbX++U69EH1tgAsSIF0uBdjk
cX8l3ydNEARRmiIWR4rNi+xXRBeESXKr5bb37ELTABn0Z4oAHzs/IV1Rs8q2Z9/iF5133+K6fhkv
bA1722WOiT9bhnRQcoOXNxOBrxFtX1TZO7idHIye7V3wZ6jR32TcWQ/aDFGBT7iuBXWiWvwh7/o9
VAQAu7O9+32Hek1RPgjLkV1wy/+gNwcfm2zwYSbIZXVa5mzX4xHriyhiwBY9Yrb/cEqQE1iB4/L+
Po09EBi6p6DG/Flziz6ovfUN/6ZslYD0uKAEmGmauYYo3pWKzvfeiZuRMde+SJf+9E6M6SoEVnqA
jgTy6MuCpkUTJ0rGHZn+F73e/gxPTXgktEuKxmTTAOrZ02hPh0WH/6vPs1qwFfEGzzqOdV/sIy02
dJehtAQbtd+U35mSyqhrnXWGAxumWKuen3WyOyn+4Z0UpkBX6q61nozAYht6sfqRHwC9szhhayLF
YjNlYkr8oHLzfZ36XOSifvsJ40STZHULeKbYbPGHFyEq6Gs9ybjnlhtu2X6LpqZDFu04hziYThtD
Oj5zgyz9OO0ps/r1HaMu57ZuIeEVszPjJeJSb2JP43hsnWCTi28K0CD8jeeTL1gKKV6+upAIlX2r
gFIqXV8VqQzvRXNv7/fuGoH/Ky6zwGAPBS2TWRpIQMEUAungph1/bMfv27XjpuBCtsog25LLvhFl
CqyzTNmd3CLt8uodmWmnbc6NruGtJbvwz5wuAtV81qNDv8jc9Y0wZ/QqdYogqd8G1WlIX3TztbKJ
bEGtImXbGBmSv6kpRFd7PGeQrsaQcmHkPZiUcO6EtPhpM1ff/x11Q/8TSd/i253salzElC+RZmbv
GAX9d9JE5I5bDg1j8AiCng23OvgB7QSX50QGp561g3UNlArGwU3bRp3nuk+O/PAlFQGn/ea47TK/
deJCfFpm70kb9zvOCtXWwHrkgnkm4k4zCeIEtnopOKj6YN6C4tlCU2ZFxPzifqb2Sp691cUgrMA2
jihXj9h02Q5ZmjIhLJcpH5u5YfOwC/GlzUHbaW4l+E2zdQKN4UXnigIe06nJQdNRagOKqwbwN7Dl
8pxciRl3libvGMTi/vHHvaU1YxCHgJxxNWm2+V8vnMlzltzU9QVC6zOrASmJAAPpTT790U2su6NQ
6zM3ec3h2bLot1two3Dt5uYIIYlc3EqjniPAzi2aA+IJwSy9qit+ItrkQEzJWF8VMQICh6Ah9Eet
caWjlWGAHCyPxINGmgqAM7ZeHVqCxv3kJ98/mXfoa4mLu0eX3Lrocq83UG8IAkAkd2wft2P/IhZ0
MH7EVBBAsRlMQPEpxwrc7gGKAIgLZ6mhlSIgQUhPTSSjnzgkqbbNCecSaVQJ1f3Y2Whps59MaG77
7UjA3+zkIlhCFMcPJkqSrHa0dDl/HFcy5jOugxbbCazqT8qqPMlPVV9cxNe1xhl6e4WwO2Csy5TK
/BlnlMBfpJcl2FGxkM9booaXiaPWLxv10gAyB93yLz3ZO8DrGL5uhu2fQYoj+yegS1zwizBUlQiK
PxQacxFXYEnpfFzMNMACA8VFeFbFGsNNU4wjlLZ4lhd0Ws3Z1NxsCbv/EbcujDZbaOaMDQ1oQwKx
epkx3sDLIKymMaOYkdqEcyKTtUvMOlKT4SCeQ2w5qDHHw0vZaJnBKaSN3x/G1+AQXOj4OKDcDDLu
fkiKROyKYy1kjnrwKurtNjCryVMyLOQUHeQAP4sP/CWbBfvRfwbdDDgOFxCBGDmDJwf4ef3V7Hbl
2fXQgs+RA5/iLWtDLJhGQGY+N8OfDGfgjFt74ECWE71DkN7JF9u7QQpwRdNYSsXtj/BH7XOrrR1L
ner+jJBxZwsuCAHx7oA2mnsYu691bX6knJ31enVbYmp0a1ZYyXHt+Xe/8rn5uGjAlEe5Az6o9KQe
j2RwU/CnOWLq0Fy9b6WicPjDutj5SMMRujz7mytS03Qs92JDK0q2rUKd5HrNtx/bSyBa5TStwhTA
/B7lrOMqaibvpOdRJ/UuDif1khoqjFszUM7z+1sDgW32G+iAbWexmZZFoi4Ulv4QZ/QfA/7YhbK4
7p4XVHmVA9jPFZ8K+JPM1KcvAMCIdCMMP8m06mpIbGctJA6gY51JrDxgz09rR77L1CQmqzdvkK8e
49x3Hw0nrYccalFEyblrQLAivNQ5LIc/0OHGVb0IATxURW5UMZ7OD+8HCRnIKHDZ7JnTuN9apBA6
huGny1i+ypDPM4TOT4xfmJsUJUNSproi64Ba6MT7QfoyTvdUxeffx0h2Zh/tDciSCaN5KL5+4gON
DvRa7AI3RHPae4ybc032Fl39Q/ppldEdKu2LnUStn+Vc5vP1T6Yvu7QmGKiRoK7egarVklQh3wK0
YHuisJzCN6bKA8elRMfUbqD3OdcooExRYfE56gJfsi+CSJpihmqNB4Qk87dN94B0b6sYZPAyzNXn
C59HOey0li44DOBrVys9XFDv8NNO2XzST034+G0pwgsX/vTLCFk69ZNRU4ZnKzrc/axHHpbkPW4J
+3W2nkQouvIFjJ8UJZNSJtHrf/yQ2aFQzfKi8gS7/mtFa93+ptrdaQKuEyrXPIpBvelsnDd4tTSS
SMIhB3pShE+NqCtwtk6+9/ZfzGnTjWha3TY3WzXFCMQPYZy4KI1JCPYLmrzhdgOK/BbIyxE+O20u
aUg9+NHTvG14ytWqyJQvXyCJVoy893TKOqoNe2hyEolQkiqAGBTMrD8HL3TWB5NZ1ZJjISbizlrF
bg/IMOhRWBTg0LQ0IY1AWEftDgKOGI7GDlwqrjwsnrifJCw+SALbZn3qyBJboM3B5tKPX2MsAGKw
uG0T9cr0YIvLGTGhBRIrfmQaxtsTKFSIGqvmPPqzjByiYEYVgARV03OiSftGtFAIMJz4FIbkFvjd
ulNPxFVnecNiLBTjsr5Qo+EOxBPVMW+7rAeoEVZ+/JC6z2Vf/pGkmTvBS8RkQrUUKtNO5mwBOUy8
b5/ZxyikHoKYoqoWNwfMtfGMjcZpSKVoScBanaLRZsalr5ZZ6mYz8YcDiPKPf/8945zhNzpXjQhG
NU3qxMjIfXifUeM21sX7pfZ4OMIDnKd6Gjxm3ePNwveJKVO+CBmv12MMX5j0ltauZId3tZ+VU+xI
OWkYX1GHTv/GkE0ZXE98U8mXS/Q72SRSGwqtuhyNCm15jbZjNFeMe5dAqhItk5UusakRbfo5zGZz
2HAW7y1FdS+TrKwjoJG3v66xdbjcNwmCwWkG+zrfrG1MDMIqrv7Xkiuu64VKJoY644PsVXRt6zOl
zkL/KLbT9IvnKIpT7B+BcCbm7V0qfaRRxGWwLpFFlN39Nr0epnuOjNpvbLearHJjo7BruXRwKXXz
q1Mo9+XXfeQr1Gp2Gz5nGESM4Z70rsZhMgfJbdB1l2Tco5KeFlN1/CoX8hAp/udIRy+0YFwaQPAA
PVlUa3VzrM4nOVeF39jjf3dCrwkSQBivM5Wwz+l/wT8zrb43G6ykp54ESR+syj/sg2zi+5W6QakH
i4zXt5XQ2pHdlIjtXFy0iGDdYPOnDUXtZ7Inj0xAI4zMODurW9PDr+K7L0WgHmB8nBMZS5BKa879
02TomLzFYgda1nVwJktDj6XACBw/lXasRpf6PAtA8rPfkkVjwSlCs4Kx8jfLT4yfuAtLUUrmYas/
n9G64AuAlEknrTj9J7A9xC31n0bqZoTM4gvtU3X8DwPHRJ5AxU6/90srDFFm0Ek6OVp904DHvUhL
sVfQTCUMIHFqOdubC/roYu97zLmmcriBJyUfWyTvajGCDPZaEhsbkD425b90mMBe330Bo507O/4q
rgEGXS0q/NASFLb8oz9apMiNO1iy3vS8qYZCcdW+Fmu9+USmwbUHGq+klz8rSyZ/Cg2dIfXKXR0z
aPS3VchzsKkfkSdrDbhmvdnyZ46Tjaf6VGLzTQKS2A2VdAXt8cEtjvdby7P+UdvR7dBFN6mA33mN
o90nKPFwWlmgzpxSeVOU+hdmacbLYpouSNd9U1EueclUvbc4MKcwu4iJ1e6qKUccr4qSeTy1vHi1
cD2zRXMcl/KQANiWVBBcaOYm+R7lohVCYbXLOUL+ETn5ogX/IcHSHev/IiD7cZ92WSVwYcH+w9P/
k7jTDvgMsqu8oXxUPSG+CwEmJ7vqfNrAd6Vu7D9PQAU0blFXINefiTereiMihAbSyCcCvQF+ODGg
1FdMhsq3gREwASz5bibZFcg7vV5sZHbty46O2af8o5IRXV2fZ/hfQNvc/SCG/4s/wuoYm8LXFLr0
qvUh1GZndIK5ralmnuUgvxzlpyf0HszuXURVQpE2FbvxlB7NRM9OfbwosjQr6GE8cfdQdBTKhkw3
O6Nsk27xBOuCYnv5usGGOLURitMpx3fiZWNn/ONBtPw2hsM8f404K/HiQs+PlVFaBDPoP9Z3nLI8
n0axX2Ww5IZxfg5RfTvRlZb3UzkCmfXkzJvih1eBUdytueDry7Yezt0DaKhKM536zBcxYDGO7v5p
rsrcY5lkB7tEUNleHq7c1xSuVXPod0q+sZHFWWPg7Cmo/2//7XEWBhmSPZYSpxU9J6CACjiSWEuL
iZCyiLtPcPAapGZvho5THsfCx5GtE3aN/whHOeo1JoWcHOlwQoSJ/Hp5JaYC6y1jMSzpdY/rFzf2
q9jprhDv5fU0wYQLn/fX8iI5PUtvV1bYyr0hjC7CXKI6eGToEMMkP7jrdduIkoZo/W/H8E5hMZOX
0vufgbBFtkK7R9msztduYca6MZB8Kfg2O1EkMd/8+f8jJgK+Wkn4u6fUCTbSc9o3hCiuqw1NWyJu
jpSe2xMwLodOAJQGlcoZrTdAZuMok4YoNjofW/rDBnryURpa1AmkJZg7NPP07M9UA2c9aKT1zCJE
HkYwe9Nixa6+12ug2dBzN8rTWmwws+UyGYe0zfAlLAUzV3nYphM/V1x5j+NimDhYH75VyrpwqccZ
7XCEkqhdSV/Apuermx5TyPg8JIkkYO/CxwdIWacYjyINggtLeg2Zi4eaP/8y6FYq3c2z7UX+y4zu
Gw9P3atd5ecjt5KW3Csg0BaJnW7rQI69KUix1aQGlIvEVZ+wN7LrEyj6MxSxPzVq4n/1jA/Nfsf1
vnKFebUzwv0MWjKm79PrKXs4bvuxeYHxRgSzMr6N9I8CwqXeaVNzIGNzRQ0Dpu7jKEOBZRv1WkNG
sVhV1VD4rinbYPJT2rxAqY9URqVyvWxzV6RHIPXAEAF7xTgdjAnslAVaYIL/Cn8riAJwRX9xZ+pC
IWzZw3S5XqCOaLgzzENaGK4m0SfIATBNZ7pvGz7zGaF3/1JEJjWadxwXM6lh9x7uDOGekE/bduuW
EAoM81d0R5FvbfcQ1OinudlPY805dArdKzdce3TMbXouE8CjwhJ0LQiRPH6q8Ko75EiAzXJe4Iut
RPy+pQV48yLs2tXFeaxFedLXv0wn0Co7dTu8k/2iPpumHJWSpF9GNKlw0kLxoqEOnPuG+fwipVm1
QCJgat2f8PSwYB3/dFl/tmA6zPuywkUlA/3r03lN3S/j0RmL6UJsb31rQIJu+mIw9icG1iOUEVE0
fNbqF9Qdli/WpOJ2exXcbPiIjQ20Q98y9ENUZdi7tn6ktACVCLL+MGIpv+VMTa94pDq0mPUBxUQH
biztGBpg41C90QRI1sisYomn/tS+7yo2dRSyOhCypNC8Ji1bfJaoL/1sTX27O2ULjSRCkWDYtNu1
+nyKXlkbK8xPN5zdBpxdCemTJb9r4ubhDIW0/VG75TG17xL124Za992JJ59fq4KkV9A4qDfp0z0c
JVO/APhqbN7EAvDLK1j2wOIAWUqDYwPIi49x58uO29DcTfoqxpCq7yWRqzOhlAUMKcDxGhhO2Pfe
4N/LGqQW4WzBa9lXyeJZKxUdv0A2gBNHPIWJWYjijKDMr6Cl+2N4JmMmgFxOcLaq5TDJ2u2PaXkV
6Pc7g2VL7go8J8FNWhyzoJ9H4D47ukIEwyJyJcfiBOb3Gdonul/JvXpQ8+HSmex1he3POISrEBY/
0MSFQtYw4V+3JAtrYRLKi0jBklo11RSopE+OGuiVsABtbpJJVdx/ok8TOxYQ/XvQ/nyP7/xQGW2r
rM++iglQ8zfB6fFTwgSDPlRdKzStyzrMyyyDQX7ZHFG9/46TMsdgBewkMndedCDrKZtpK9LFPBzO
Lw9/bB0EI3vUSQ+jwd53r11HtgofcpPGSc2sNZPO4pp8XM8Yje/n9TUgbflMglfTHXnEGdTvEBRo
dxhzkMs4ctKIWNgn15iiKsOzG0VZfKCQVOScUfuNUX5Z3/TziV3L3WOAerVCwNDkNDuF1MprApY/
TkCNw/Qk2gqjMy953tgh9a36FpPPH0HVoUq8+liko6802K2JJtCLKhR6BuFWxbhW7NXCY1gbmMQK
aIH9TP2Xrj42vixf70tDZ5gCxsiKRjlaHGgAw29HGvBndH1vX2qizw0/c0dAK0Rm3wkEhwnDxZOK
x9zxR5R9nZ9YYuYZi0uhsUbDecQG6sFS+p30ytG37PCOluwHrpWaE4ymzwFqheQAFjHVJOxylKB5
sTYVtWnXM79q9VY4UfHwsSFZQu7yKVqdWsbXbiS1J70qELHXABZp/wdwlt4ytGLkoXZJk6ltDp+O
vN4oY8mXif4whbPsfcOW6lWGQHIbhfAp4eiOeS9cIWCnTER4WekwUHvB4Dh7dbxOCCsQty4MTG+F
OvPUkRsjjv3hiq78BYdwYbcEbAqtsSfkVlwfdRP+U/qqg7WEkG87sO4KyQUMyhccaUU/sG41eeSB
Eg9Q4Vg0LmD0DAyzGKJ3eiPD6My19BMBwmnc3DD1gZTNOyWib/sm0Vr9soxc7Fp8xe9FFc5PctBG
aEgzpxsV+ZaWRxUHgonq5nkYf+YZOtxQ4P0ivX3bMmuszXHxdUrIPbRdsz+eaAakk91oBWCmVdLZ
pS7d7Lg2AXxEGliYjV9k+s+Z4BHMJxuM8fxccEYLz57lMeVDC1ZIfMpmTZ+UKICNTygDy8Wb+eTF
e/mrgfDs6ly/H4GZ1SRD+9ncXec8xZgZMKuPWxDLTLVtqoc8kdq6CcCvLrbNtMMpvNSwogM0crpu
Uvza/ou2xR+bo6o7es6bD0zwxlljoKqgc0cYtnoKk1eUX+p5ULJuLb9qc6ICasvr4zAclMIG4utj
//FMLinrgxFWGZTVHnhr6iqxTgIl2Tg+Z19Z4DWtlNmTDy7GmasNXFCMaFyDCqWfZI6m/BDD5xsx
wPqnK0htod2GWPelQBNjXqqtRsGwKo0xHufF0fJFwLpmnaO0FlS+hyhxzLD9UQZ4RNaY8A+7p1Iy
hJdGr5Jo7D5FLkfLkZSXvtGRT1ss8zT5F8ff8aLssNMHZYMqFbG8GNVbaNLvRWpCoyz9LJHtT/q8
YZvP22qmA5w9MYnNW0nHgKMUXXVwIB0RCFc9uokVRxFV13IhG6IBaA52ugDISH5tHmXBjRbOIurf
l0+zD4Rx2BsZQfhAksTE3EuPJeR8LkzpavjqlIQ6J7MaR9JVYNHmHic4DPInm9x9uzhVuIVJ0eKV
WBzmSghgBKZvgjfUuDWColry2Dl8Vkl4kNs0jBTGhISiikwSeBmPFNWg59Xnv2g2ukLPmjPoxoH6
OPEsWUVCcQoDtC4dAW27rIZubLa5PCsoBRNMHqoVyMdEM5vx8sriszLF9Bjo31WV74roJd1lbNPP
J3WZlx+Xmrnknhriyxt38cwbm7fRT6CUxi4RoLIBuQtZV6npzxUl+zxN0hKDZ6XSVawysWpqlpDu
EOPz3m/fhG1j88RKRpVbWFEuLZ634IYgGYE+AAINrVKSN/VSGNaKcNkH05DwggU5HoXdYH7YG0xj
W78T0tjSIHJhXY7VonkVS6zucUGsRy67NerWWJmqrofrD1suSH+Q06h5/5WXfWzbZYKO85VLuu43
dnbjNgdfcRRg6YuVhQx4umET7udfnzk8vr3+1acWcE2YwzgX7zJZLNu/g3fuDMsW2anRpB8hT41P
UtCVVVL61AwSvBBm4O5jGG1+TgXDRKJkESZ8W+R1uQeSPi6HLB6VQ2wb94+BjfmwuFbQ+8nSBP6q
iTGJhWF5LT3RdUOQvsqtfhz7L4DFpesYB3toAT7zJBwflRUsqb3cEnCFDU0BRLabW0oNhFS1goiu
ZREuIjL/ueKqpWgn+Nn98R9kf8fDw7jkTuiauqx0cdrL2A9LL5aBnD/fTH5DxwlN1y3K7n0b1zRE
BnXbhTB/DAlh2PF5K+SPiSNYhvPZzWH8lIW0I8WMMPNO9anaVHjRwfVJw0wwuqMYXyhet0/5GZbg
FqPYWp0MvTn9eUs2siSyzk3bM09W1KlmmGG4Ei1jk9QoDR3IzDUPpj/Xc7NIgJqqgdJhyvyBP1xf
c3SCJEtE0h1VMraOzl5qDksli7OghcC3j7cZjuiU456NHCCwUKEJ3JCAM1CjaaEPYLiZqq78jhZ1
Q7O+9pD8fBfY67ogs/aMyMXhxRefLJ2AupuYuM34Ja1nfD+FWi4jmdL7mpkKEatDTFMkMBgrkL/p
gUd52WHUFZ2kA3qfugLv03fcrZR0C0OPSKseB5ebRSpt0QDVN2VT7cl+Wt/TG7UKpkkrtAN3Og/K
8jPBqLkBELqkyGN6hYBKwq2FCFpupnpQUKYqRv6znRTgTZ3NfxpEibMyvr+efmeNr1AQzhgAwYKb
NLac2nUicz4lDmo/2VzA70R6jomLblhQ1UHeBbDgKXg4fUD2jT9VeNa6Mmzc4x46ODmRvSsrYWj0
p08DzD2ieHe3hwXSjwmgGD8qoLGdun6Dh97kMaB8wvMoP52yF/7hgbwizWzxoMR4vcmhH7vHEJE6
uRzEY8tgTw0y0VjV8TV/qRjYButP4lIF1GYI1WlUjoVeQksp73uCanY/TjnZ4Fjndq6vrXRZGRQR
kyG2Q2Or2aKOGxZwqhs46sQxl5nGd2jBZMtcPT0gm3CQ0xEjHMUvN0wb2CR0dZAW+sdVWgrICC28
UgtjWilirp4y/S6C3ETpt9auc+qqRgU0BWknUQ305hxGK6DjU66zV9Ba/c5RlKYKqoM+DWgOE5Pl
08ZuU9rnflCe9MOi6+WiKyAGM/7zOEdNL4+x5MC67Ad1u4ng6QIscd4Ga4gF2fQMzEx9kFLE2Vre
7G1zYXbmeyfQBDp6r/Bvrd/DYqpeoSIn5JxaEs9xCWKElAX4ENqY5t46EHrPth846SdKAMxD1B1x
D2L+nSRkhLJ1BJPcRQ+5+VnCos+2LwgiLXv2ZLeyxQSUKKTZ/wNFOhycey9cmye1kn6HsqltRujx
x/Y2NLxA6xF3qBci32yYAZEMRCyA9HVT6ekSB++IYhOZLLo5onRmBw6Scz+d1gq1tWNe5EdbQzHx
al4kNn17PUssuIpCTeMizY5/oRh0awBegeN0Ik0kdFr/oByUKCAaOWa3tGqurLOSkMqQ26bDTYyV
5hNGv0E2EBhR/3B557tcac0bJrmNrmgSMGix0wzWbRnj/Ot4Pklae+6LI0nht/XrRZ8sGH5+6X+o
Lm7G1pRakxgWjs+wMYJX+smHABduv4G2bZmYHo8VVTJHz/wT/JcTbJnKO0xtqoIaX7eQQr1/PuNe
o2ybnQrzrDgc1fEFEpr1LNg+7O2p14B/tBYUseP23xb2reJzE0/Y1oPfbNXGzLXFK4anN101z5Kw
zoXz9lLvFQX7IbEi+4taLg8vZCfJ1fsFfde2fYnq77bYkal1lMCgpcsuGRf7u8LhLSDy7N9tddR4
y0HNmbl14/uFE3LfNt0eyXznPGucMplbUCOHpbmlHE/O/muAfmIjptRBpHbEoXf+N9JZlnuvN5HC
rQAe3Gw3AzxlpbxTwBRnTd49qEq9JzfLqcVFKQFqCANSrmvqLjW2hbM24uGds2yCfhbFnDrAQ3zZ
IAG/hC8099u+18b5hVWbRKsoztN8fO2ER4qnvI2CMX2zKccfO2D2Zr7RmeEaN2NIMzeGGlYCRX1R
YEGQvbPXtxNAtWKyI9MmIUenghnWUwew+ZMuNQXt4FlG/PGV6/QGeJhk5hWFFEGxVPHunqohbsu0
bI7/Rjw06TfpB5R1HIURgerC1IyExr0rYyKayYLp3KsWI3uFmcCIoJaOm84/F686mrDMFei27jxp
eKF8zx7dZPVlm1e1I9rODVmRq4+gMX8fYCneKOiL3SYNfwehpsx8C3FlS4Za/L2gFFn3/Fxu06a2
6Ts5TZ7HUgbKLXY7ds5M/LaYd5rAKk6Gf6SkT8y/ub6Pjle2hS/KzdANrXN6PrcPxgTfTd++kKBL
vaVzpxHy1/4aoivdfdVt6qqvj68wdF2NzuzlQskdM8ypWAONcfwbHz5+gKcUX6JoG8YFULP4Jz2o
jExDkHV/GtxCWgY+I+OgmvkwipR3nzd29M2xoZUD8acI867ydzx46LaO90CiR9nQA6vPtpRa5sy7
O9Demp5+bEvRs/zmXMk01z4+yijpI0xIQCo38RJVa+vuWpOn616F25+gqXyh9d3wKfG9J2qR2hVH
6d6vl9zZQMU8ZLePifLqW2oYLd/z0dXGRGg5j0URoRWIMXTuMAqq1rZG8Dq8ntsKV4W9ifumvtgd
KarIGP9r+yYMY/B4Fr9b5NJaN2cpYEij3xQiz8Pu4hXl+4H2lE65HI7mXgFe2ofsmEMKxXCKgcCu
SV5Ko5QP0ebY7fXHG5ud+aSCvw4TjEmNmQtJNwxqNg1ZO77JXaFEgewUhDC0GEOxjwkssFGn6H3w
UELtIN9O0NRSmcSNhQhXT88oghOBhq8Y8x/2wVrWCrArBeV8YVV/CW71hYTfghMC8rRXchmIO6N8
ZmGH5Ts35azK7EOLOUhcjXTAngaDBPhe7A5IEeUIqE135RW84zhe6PIc3ofUzpYNmKrn+uFAM+13
tXCLcZmfp7uTBYzsp8kNpuLF3KogL4gEjAnU67BKaZuxdHhD0/PBWhLy0AZdpBhXrdqiN8UDRB9P
oN+K4WyArnKVw4zKDnAujDKVu5yzNK5aAow22AyvXYuA7MwQSgev1O5hIh+rzNK1u/eQ0/cfl0Gw
7rZjeD1unc0NejiQOzOCQBEgBX7f0MoGKFADxRHl6ms0ag4O1Fn1t/QGnIPUlnzgJG3Bo+5xPOra
FAxaypLTYFqnSuK/SPHE8C0e5gA/O93X7muhXsNWzwLiXzSNgGF8X8r40o0Kbb3/du1efCa7PVVy
xjz9b5CX1/QgCIc03zCmvyeHTjpbvIruXd7OC0fswHsmS/QvSOAQ9Yzt3pHDGLP27rcTYwcJ2l8a
c7qm9Q8t668E5/axVfl38nObVTaj514J17InplWv1fs9x7fSkCIpS554Go9GgTHFVotaMJ+oInrf
/ocYFP/Ime4hP3eIf5ylktKEoggSQEJFeCTUszkGLRLzCdXWDhOAkh69k3ViJQKvq8oqAUj8cub0
FsRP3NKKI5Kj0kI6GaqbubD7qfbFHuxr0DO5dYod9qfi5nG5AUUTDWoHg7vsq+iCjxNQUkCtbo4N
UBgXpxHnRJfGH7VfqPxGR7kVjRd0ClilYbEym1tg3RMPXI72yOyQi5++9NIxC8QMPwOj730yz5/6
5jg9mn4UHDJqtUFicvDLfPH7+KJztHOB43yxIb291jGUTLK8LHtcr4Qfwi6vat6uwztpVeXJowRp
zUs8Vb8waOMtQL/EmPls/ron5LR4uLUbPcfWZViEv5vHHk5ymH3S6jo1TypGxfauJ3PwV/lPHHoE
lpIte5h//U1L7nT3Ob1x9Y/0djlGYiLnlvsatWaV5IfF/v3kXGjovqmWfomTZam1DEqQpn2tOjSA
EmuB5xxYpznmSR/be7eg7/kDQPGOUb7r/6IWLnuFnzRwZOCIeL9uAce70Tsvkq3TeDUeLcHjLQGm
OHzst51j//P4PChvGoPh/RUFO/IdxC2QqVTxINJj5g06dXoK3T11YYLK1mt6Pt4zIvOfJy5MjmKw
l7wZ/tIMog+FHNs6Bx483DLKVbjmYEU7+TqqcFDDeDHMc0agRE2WPxSdbj6lEm/GpV8fgozzJ4aI
Csh/xwOCxpBv9jIe8S36i5MNHJ+zvM+iXIKVtdCGizs7ec+OE46uVPCOYHrUJOE7giF3KiVnMQxw
xlyQQazJz/8SY/G615Vyj4lkQC6mmUTiiPGwRteJ4FzFhd+MVtkOkctcGE2PpEX2uoOtS7AQ4Jx5
FTQBfHaoMYlYXLruKEqAD2zviNL4WMv3TkD9n4Na90bywR8Y8BTYmLaS7eiTckQyhSSCMlqtK7aM
F4Q5ORs3GYgYWX96+2ZOfweockIarchU1OvhyMyHC32Pk5nRcPJj65r35EN2cnIzhy+HzPsn+NUG
thu3i2/02XpHt1cCWMV4IOLdunlWm61TMSupyuSddNdp/X3yCdv0zwzrJ5pSD/QMd4oreazFmxRx
NzqMHcNuGi8xNZOm99QKWlqygQc6wryl3PiGlpGrITSThQCwyVRaXnxPvTpWiyoeBd13J4ScvDU+
XvyVi4GVQLUymYmVBYG8Cy00Adf8AUjALXwJJIDofxllz9z687TVVkkxvKFPcAryitbKruauJp3L
EPlLX5Goj4ESNbQQqzhpBjIowIza6HcM/i+zGNyX78af4zieUoqSZ+JyppFZnB04bUTFbtvLPTHe
tZWtfPlzx56YvvMuvAayEnrecSD5FucDNDaZ045+XrAH9WXIKFnDybcogSIg+ScxSQuGsfgXbX4B
P2ycwajVURpDjEF1bfzKk7E1f12DorvOoMvOavxbbwMehdfztQgLPTGyKoThKLe8Qk/OqQU8xl9+
t3lp2ShZsVmVu7iM58rlA+rBomHySjdW5al0tkzF19zj9MtKt0Oi+zWstGyuNcjZFQUQdzS7ftib
0EXF025om0fjGk8MODR2pB1jpcqA/uoXB5II3hUjtb3BAp2X9LNFgeMxOLFzJyU8deHpuwX+imEc
My/D5RmuXk9QGt30V6QotWzly3HqYv9QfX14e8f9M3qQF7dKDjDs87+An6iAq5I5O/5/ZPBtRAyx
p7DIDHj4dz5N0kTZ47l7KSRcQnbQjWXcxUE68Xrtm49Q865e7zY0MF50GZH17Y27vW2LXshyhphL
BnDbPRgMDq/D3hoTgdGl63IADhzHndYPqOoVuSuVVHTAgVEEQ2wWlLsmEsTc+nzscHjxeE5Eo0ac
KEg22y1dmxZ8TcDiny3bH5YS89HiW2gTEgibk2x+O8/pQ1c2+eQg6yUHIaRoIPi8WMSuAqcfR8qD
l+QtgwFbT4td11AoC90Vp8DalnK7dy2SaxNY2ufO/Go2EbZO2tGejlDCmVopRlzgJHGhpXCs2IIx
HZe8wFc0qYvxlhP9+nd7LicoJRCE0XUyK5i/m7l1wL/OcTDFIv4Xpl1T2Zr4KSOk5xdFyUp30lS8
zz6xLFysy49PuQO3YLW/8XEECokLWD/iA+zJEB7+AieiuBeqgA8hkiJIDjuUg0P7LVcnFhfrPj+F
xhq5T0TbM3Jw2fQwSpRWjRWG70TIMPIvaI0sBsIoX2C7ggb1E7XUesOBZ9+7Tk/mjGTNa3hbxYkG
OtpcQly3AOyH8nU1pXrYuzfP0YX4UC+tWI6vREALZPRo5kDbT9JDb3TJu5XunvddyFoLM0Jpgd2t
5xYgE+bJy6FRL0zd4D79++P+0xegLINfalXUOJrskbDA2mgzbzFo+epwwQvFn2l1AekmAOG60ew5
kmbfwX2Fv5++tbKd9ubQsKzcATNPmXho4vR8FmA0r9cS2n0PoCIs0xhhDoy/9XrpmP/7VE5s/s5a
DKW619zqi2OEoi+wvHDBhUv8sXFHPWV8/FyKvvIw63tsDMlWShBLYUggZQYON9Ymc1YSZFP5fnfX
xHgfH4b6A2Yfs3e58cUm4ik9Xg8cdI9l/6PsCHdF8G2x48quAuy2J46bEQCnwnAZz+MrOODMGa+v
ByUBNz7TJIxVVMh+F0zWkGuapoUPMoeWFrXO4JOnu8s+1cMeIIU7ZJ9buz4lY1ih0479yxi4E7TF
dJ9TTMcAfK6gpqmiz4Xe7BIqKdcZm/87nt3h3Efiv6RniwdcvEy2nbG/XWvMk8fCd6oTb1I9aeDm
TzTxoo8eo2nHwTXmka/VFcFauOaXcVsxhE29P1JMkamN8ErjQhfUUYIwPvBKYI2BT/AvppzjImOu
aJoMlB1F2uUdCQvrTbbX5WOmABo8XYsIRhOphGFMIrYd5r9d9v3Cz/9z38sNWZpSMeox0pr3+j2e
2YLTtkQvuIhzQla6Dhz3Mx1XY/Bs4dliNmZtQagvRmgwQJdyBYB+gmP8/U5aNLQl1/HPjJ1amXeQ
jaPzIJFtJ8C+adpCmJ7bcQh+B9k62wN+PQnQhtG0M1TGGZge/3r++fvzS8O7bzVyZJp3fW9tpnIR
wqcrYLYGQM3U32gVjBTdyOHptNG7Qwcs9NAdJphxjJlGWS/gC08po3k57dfBTo2nZJFuNPL7gFLE
eeR1zdx1AObRTxrEvs8Es5AFeE3lAXMXi5yP8QMMPGTE3HAsTWgmQpHkN8pElRGs6yCkwFyH/yN0
F2gdQh8YVXfQ6I1iKjWTxsm085qY59muvRuK8OTLJJpEkrmD641EaSwmISvnZq7BcDAji7HqKhRy
iKpKJ6P3K0m7bwTKP9APTVzGSPBrKF5gz7XIej1J/4hLNjYF4msx6TJuiHUrtmKixs+uJcjAxkRE
q+v02glVKto0HvrBHJls1GMQGqbAhUruQEqZvEmqVgtVJJhAXbS2JtPBUQYBEWaGyR4KKBnVy0Er
jAd170HWNEfsVs/buyhfU75Ic8fzZ+JahVeFBl3lsti2E3q08i8rnvHmpa701Apqd7Teulz1NtwR
Eu55bJ5PAl2ssgH9+rBOtcxBsZFs6PPGVq+Bfy5qWHu2PENunshoMSisYbYgVcULzYNQpxEYav/4
Nff1iZeKc5L8rc45wzd/fkzaXuD4J1oE0zcrPGM2mpMLA7f35BbWMboogQSRFb7Ov9KG5lqKO8QE
r5HJ7qkfwawHPrCyf5MpZHnSmR2xBewCyjN5SGqGk5UojRMPXBaqNuakbVn9m9zNbCV+KnMluaxY
6yFByEb1MQadluHBqiMxNPlBXT1WEMTkuTbB1zD/DVRM2QswRu5y3fZgYsc4GEFDl1gf1pQy9pn8
2/9gJuiKqBiwatizOJBt6d3EYSjsq2Qk6Kxcjm+S3/+cK0q8sGtRacY+h50g26RbiWqAKJDbtNZm
VFu4oxwRIEb4H2ub/EN46Ejf6xadD5EyqcYmPWo+4HRyNVUpS1TYcNHFLo6lsgEMExkmDaM9jwRa
sMVIYIjB0io3g3rGCg7eDTJLTHkaMckMibCqq9eLV7atqNfaQc/ZZSsqmruNUWXnKD5Wwv25SVZi
Wk2EfdTlY8w9ZhY939dnlFKIy5mfYXaPW3HJ4v4bMiMA7+LIGXi0bExZv/EmRWI2Pp743fDjKBVS
WX5QSXg3YPpymN3eO2pTlzF4NSpQppF+Geo/nuq4XPP0Uh1RMwvjh6bOwc0zpwslQfZERzVVNZ71
IlVEZ4JIRN5i7ljlgsyL1nNg9U5a3SIZirqGHfSBA6X7OC7aRehIEPbIXSJa17lQKgV+cG9BxHVr
31uThLABO544z8vYXKpsbOxr4DSF/E4ZHlzTgPfzgXgtvSBigCrGudHsLo4Yn8a5FWySixKxRqA5
02xFM+afy/KzYfqkLYQZF3K8V2Pyqkl6kVRhLXQOlEN/uBusybkmtIRlBP2+sTk3W6C41Lkgutci
niK8VdnkjH22QAlPxW6ljghQgHDLMfxHYPKe909oWed0ZRkuplndQdMN7M4Tfa7MqLcrgVFEVt9Q
iRfjceTZ3suJEwxdx3sI8VWoZsGf6Y/uR5HLFKxJaHGL36z/ehjStPRW0p9gu40ACXAMxjoICG9m
Q+0MBn2JCdsaWFs7w7q30sRmnyFEEm75VOOQ45WB/rx2wlxtfJoXdqQfqUSMdASPVme6P3GOZieJ
ZMdN2kZTzzF9g7reHgZOEmdHKITjb11RvanTXMJrfyGOv9rqdMrI02pgp0sHFiSqfYFRkrM5ua27
FGQ2UYuxge5Ge/D0UUh6CkR1l+M6LCgPw+ONqSYo3HpbEb8PUrJwxdujsoNjPddE3M9Qfr+Lu87R
4kVCmB6Yfnp28jCTgm35AH8brTM+c6aWejXPO1ELKh3QC5vqWprMsjIb6zSdh9O98c//cEmRIT71
8rkWkq4eISoPTa/bXE7xLivLtwIeanuus5cnlfu+49x6em8Dm+rzIabvJqwCrtmM0xVz92txIiVE
ggo6jc2Ri7mPnUrKtOdCeo9Xc9If6SViZEoifihEZUL8UJLL15msFf9WBfSGmJGpdV2FxAc28tE9
zc5egz0k+UpbW1xybiRVu+AWzet15k7D5uG1SYv7AK7gdOO0G4hNmQaKdfEepIQtXyWlS0OFLa1s
0uHriricxZhJH24zQ9mC1gn/d8QJA4qoh/aeTZx8rcVdAScC04b0ZKJztbymMZ480WnJ3wKVIVOd
loOhQ/mDPqi4V9YRnTxd0eF39LE3K7jzF82UMiwXQYFIXrh4EfV4VQUGzO4JbdcNHHQ/BykS/ejU
xcqYBBm4U738+kj/L/UyA4rwWsrQRL8ml2NGpPmfLjE66a1o5/AChgfhO4lmKqWkrcNJE2kiUsr1
ob5GyEwPR+pnjvXW6a9lXDg9Mi3Ie45MoMQ0ylJe2ioenKoZsE0BlAv9VVxKyYjHS2/cj5wU2EPb
v4W5+UEBq5wI5PigoVqGcXS6g0jsdmE08us4U0MbF32E6q+s1P1TNdkV4F1460JmJH1O/wdoplCZ
g+fVbL0aJAvcmmyErK3WMoeroIzw2XvNbcKjT3NCVmW/lQ2F4xKNHDdAtOYl3etEJ+9ckRhnQHYE
tPlSjDZjNHY94nXXIekeoNRabWuWFz71Rha5H4Jo3bQqoc0YtlVBk+w8Av6h9GNtZd66F4dOKcV4
riEkqYEEMclqvEDIj24/7uKvD0AGQoFGaxB2/ETqGnx16FDO4PRX8yAh2tSLLA97Z+aM8PYYHedB
RdXWkay/UnmMV83cFnGmp5FXpHbpWFxxlwGXt8bXm7KG0bvhUBlg6jwrn73Gmxfws9+gbQ7LHAN7
a6tFo9xzjtloO+Ulp2eOTkgZ6vpnsQGVt1FIQk3NmzeV9vYgmYLv3BSgrTh8/nO8l3mS2CRXa70W
gkYe82dxOf+j2QO+F1q9+CN4LTw0YGPmh2+KQyYGKzkDTJiOOpak93t02bltCzxvPmmI5VfS+8tn
Pr2WqF+D+MngdwosTET+17tEMfy0cR/Fjasz/Mc+yqFha348irZCYwtriPaZgJ25kGZUOm7mNf5+
bf/DMU8dQmZ7ZmGpIqud8cjqtUtMO+WPyYzkAAXwiANU5y6jGFbxnhGzDDoVVNO7Cm3hKRJsXJsX
U6Fsojx6SBA9UEF97dWXaDX9yRNsKts1KThR8y1BRVG0bJj6T/shPHctdGJ/7ODY2AtBHdgttp4A
7F+yW5S/mWLwpF6mm4aQ6cbDXQxqefWXjYMvhUYh8eFbO3zQPXJQzRoIopqkNz3ao3KIDBywZFpa
S6OrLimIBupubmjVwZJD/zfpC43IfHBMX3Xfzfb++USixgKAhuPnuSPpJXP8hSfmAK45SCTLCtUp
KBPuJPWzGLmuWx/NHVp2wNCwNTOSJt9dh4ug4jun4s/1UHn5SXNfJZfAQqzTdf9PYYmsA2KBuTOv
J8J3OvkV6b8b+GtKUd4lUQKFah8YKaR1DygCs7WfUydrVTGWwpL5klmeCfRs4XhkjAbX/pzjsNMj
zdHs92e9hdlBorrgj0m94erUdeefziPxHgSu1iT0pHZdUJQBIEqUylcOzGXTZrNICGgCx1kEYn94
HyhL70A9Y0MY47Ra4+B/W+ke2mh4xQclklJMcF+MaJjnD9xWbvcd0l3jTXZi1ueujKnRj479n3gj
yY8PUMguV9DmJHP12aSBvB184aB/5dtsMICb15ByzwJGJld/FEHkkeOtZInfQ9s0dH0A+bx9KSfo
hVn1bK6hhuxRsJ3/Ud7il7KuRGVpkwH/pAN8VRbbyesq9SI+2NoVH5jvfuE8taOPjY/di7gEdbOb
5raXrqVIaECkZ08Qi7nlZb+yn3dbjhwNwB3dFeCw1BEZPgfUbLXQSNObZTWIICrH+Hfy+6Ktqo/H
grqTfhK9GrmYGG2jAOd0iDIR/F8OrfJxYh4tO9nzL/PbXj90SQyEN5W92tURie9MbLSVsweOD9iq
M4NvX80pJ47r0HMCLxnvFVQoj7CRo45oUDTflE/Fo96Zxd1aVXI/RTlFEvbC4HNo3d+l0qfa83Fx
YBN+dsoYMS2TibbuqE/mM2Mkq2kKJ8ESs+pk3DSCCmpvyPrSOD55xYwoRKUxZSZkYnbatHbusV0B
RGmUPuSjFUzOQ7OhbIyVLpjfTRN8DNsEr+zIM5mPA5j8Q67kE9Ek8NzNXrm14Jsh6jE82oB11vir
O3WP9DO3lQf925zzuQgnFEbhb6BphM/xAGkDrSvT+5wLfJtasfx2y4LTQStnX9OeA+V8OGGvV5Lv
TxU/4966JyutE4hDykshqBsR1EIqGuUw3GTvHbj+mVFsWj6Wx8caBZ5Z4abxu1XSyu++rUtDQ/lC
93x+hpUMoAgzXzLK4kFUKVa3k9SYuOPrbPJ5+O/pMysyvT2HZBmnDl4KTRCFWyjheSOQ8/EOcYpz
B8l3WBrWghmoK1558YG0Z5Vg2dnbGg0ZlKmjtPRgkf/rj0y92q+NAV10gMDXT0Ns4YIevPcrL8YA
sRMlAmcXNp9iaGstVUCrRajOrXVIPl14pZWGpsKhI7Ukjk6JkST57IHMhfdaFew1IKXhatvskqlK
X3XvXFmnjbUfMaHjECZ0VMHgHPYRsdAVPcefDbTXOGh60VrD0xh4AYUtFMoQ/CxNguTmUfhPHko/
T1urSqrO/S0OEGJJFLvH0lV/SrtJ+HlmCR1qESYWyIrGdStA3D2Z4K8oC+V2VmABWtxpQlP0zTuD
519DcorbCPznbSaQsVbNAviigfq+rwZmYfOSVgTIE7ik4MmSFkPvC0tvOruvX2KseyB0uuOclKnJ
VqD/7TU1AyXZnCE+4APTi+Q7+bFxWVwXqRUsOH7yGphwus1+HQcHES1Ovd69tP03AqLddf0qYCh7
vMZClhT5XOCOpAxwz1UN+H62q/BCiQEJegf+DLf5ObPqB3wuFUObFDJz/S6CwYja61aE3EzZShax
7pDNq9V6byQ7VsB6TArbTw7XozMbQ7Y5hCuhOqoR9molckofk4Ulryc1fqNO7X9wc8BEXDaenyaZ
CAuqoqCONcgJqgu+e2DDOgpnR/cYTou6zLfzC8lTQh0/JdTj0ceGp2RmfyjYAh6rRpLq8985W6O9
ReUnrVXQLNTZ4bLBivNY+njQM8U+VdR55u2J2LVG2R1ZCI6zZHnbl961bJG7W6K8P13owLJ/hog7
qrUrVnuG+u8AslJ6ZvLifNnilWtsWO+uAJDos0EUVrXGoClYA3fM7AW+6Qluh2xvs1+l/bdyJ0Y8
7h0ytDdm05FN/tFvu/VZd2yIJs/CN7aiig+hJU4Cntv5GGnR31ivwjsYIOg2L37B1Q7NeJGXs9xR
bVGKhU4Sk4Y0OpBOqf1ht7lWltum4LAou3IXyTqQBMmmWc8YnlakkIZxMMKcmXwvTFnygibiZRO9
/lV2q+LBH3YqGRCWCzsuBosYquwp5ggk7mZKukuHQAkBE0ILZTAYpL26drJbVfJDKVztjjsl/Yue
cbLUvYDX+/LEI+O8C1mCbCy2Hdpmtmw67CdaVM+rwBdKmiiEd+f4YZlgf29tXrDIXA8Clrs2ckbL
m6Y6B7rmGyldzo78RyH7yRW4hrplZ1fdYa0rc7N8xHW/CRvpdRsPxdFZgb/ft5F0vw3eiLnjPDL8
paLN7tDqMJydi2ZlSbQDHUsFGJDaiTY0lGJ2i0wDfA5A6qpbejWKL/tMXhU9Ubi+GwV8LFkE1pVc
EOfnmNDYpLwGYWXp6WChBoytmjJlTkWRWLCa17SCHjwfvRrO/+vk4V+Ik18gwB2ZsxOs3O4bLwig
jq91ctYawlHUPOjlM9vmY3FSvxZ1EumqKZHEP3JKDjL8W7Z/gFdPiBmpWk+R0YuxXsjtQTWFaJKb
9dL0/GLVDPZC8QEFzkOPw3NTu1sbwTe6jEl1UMa/OXvphtNSx5lj5eMjfFzpUpSsL5J/CKfJeUQp
JCleBpkb43Lou15YGyLki+Y5xBmsEqcY5ZltVASkV1aYgmCHGmI5+rMVE22p/vlyyimO2GUt5QNi
kySu5JR69UABKRCaeEAQzoSmytk530M0MftKt5J1/7GT3ofbEfNb9I3yyVR8ZR6EFFrTnXFzHf2w
QPpNjWEpiXInv6/ogJvR6AUgmcwTc9VzwGhYuKCA4Zi8ZhiCQP2jQAp/VhuJ3adt/8o8+U2pYUbU
bLZmvg8Q+IVUTFsW0NZKK/SJQBuqO2/n8p/XkmflGLg6KdrHO/wx4HyoxX8rL95SbdddwdZ28m//
dV5mj/g62+vTJI92AQAd+1papI7VMJNt66NQnNrTMlg/rTwEQt56XtOGUkBELrm8+iec3yPcvzTK
eIDV5Ls5P2UKAM9zbu6ulY12qI8MQgWAh4GVA9BqGZzNm6kT8KMh8C6x90tQL1gU81hJsgCOZpGg
dSL9rnu0I9ujTmmy8RcMCf13oLhT6BqAimgpHlR8YtLW9GHZZEzdRIAOOpSqESsAs0BRrHWWigmB
hS+OjzctPxyMUapbMADCBwg5Zg4zI7E6yvDdk4sjZg0MbqrBMsrE/vLy4wQxyGWwTRlzG7dpwnql
QtQVtRgo8zIP7NqAh5fy8WUlBWlES1phKMk5HwFANvQ6dYoBlE3LJZz2UdlZvpTm9JfvsjT0Ii6a
lj4dt+SkE4+VTSIu5j5j158AEDR+NGGxXZ7jRMmu2VnebDgeDNjrIeCv/tFQuCigwHUhkQATRe46
/K+9y9yqDBkDe8zKVjF8nmh8OMm6hv9aWS/e+5Wmdqm/4IFKLsX1Hf4GAjpK1p+mrXzzCDHLQceM
Jkjx4qFISPWB4PDD8wkcm0tH4XCrEotW95UzkeK3pMJU/ezu1NWhlRXM+ZYwkRPflTPqlJV5rBM4
VxHsInF/0MyfBjWgjbVs4od1zoYGtmnHlPSdGzXcZdZeTJUiYxlhy5JdEZwSVKqZ53oauVGguehc
l9AfAYlvkJ7VEgX4551nTUoRjQRuDS1OhqQcVoS/aCDh880xL3lpHxj4l3laS29wiXc4OMMMAm5M
S0ZWoqP5O8rrND0WuNfcnxmrmM0H3HZyZPKdf6c4YgZ0G8pS/DbRNP4jSQJ4rSkbOPFqI5Wf8Ibc
GplTXyVX38+0Xj4UdEabboD6drp61/NEk7VSTgpIgx7L22Z6tFL15bRdZZwIoDVcD3U7ReNoz6Cm
dF8ylWEaV/eRVKAW0BTgeBn5cI1h+hsMHfqEJjpw8zAySRdJz3WOC+BKRN6Q9nBUuInqMVATplI/
0kCo6kFOiMREdm9FK3yAZqHGcttUPFGz1bNaRqZgB711ggEBu8BnQlGYQVfaHOGXE6VPSL9KVMHg
4tlUMPnOovI+5/tEpxdKdJWJIvjVlbIElZ+8t/3H73r9vuNpuRRlKW1xrm2v1U2dC2cmWvXFTsEV
hDYZGuatklTsC3dnBPErfgYinzKIFTfGsvxkXsjPruIOrikA33r/lSR2PpIKRFiycso09L8WD671
pThZfvgtAnJRS3d7mH9J6X5dccT6ubvHGZAXoa0ts4iLV+/4WMMaMV/bl+1H8zf0pxcPBMy6JGnV
MmZTSBAwoCWM4pJM7g3mt9aLbP/WLbe9i6XKL0CbdhdDKn1Fq7yRzScl8giKB7AxdzjuwCsD2sh7
fSBuZTLuGY29ryqb4TQ6x3D/nVO2ofOil/NriL/6y6dw/WHpT92lsONXGxdk5bz1XFOzMBfL1Oru
5V3Si9p7t9ycvl344GfBlODq767aFfileDUy8Kb4xtZo3yDPUUtlX0/wb6nnZQWQvmQAMgOS3yHo
XqaizSLVu4YeGxaAWxPMotuHi2NhaRb95QlpeBuNVllBldGrRPy6PIPLIJDZ7iJUR/UI4GIehKph
01MVNttKcuiYTZKddc9NQ3Pbom/oRfVU9thh2PeyUE2rvDQqHADmFWP4J4SzkvZ1uecedP5urfQl
YP1tf16sRt1Jlo9oVHIbaZ1YtOApylDNx/eSj7maZ2SoXF4dNc0CtvGCQ7qNJk2BBIjp1ZUE0UYX
kfyDENE+QdHvLKKtVUm/60UsoY46ITupKkX/eTbRS/4mdQpGFxTfV7ljKWUorb1O2QcGrU/Yvr3w
75yK84oxMQ3/r7DxYmbhyE1m4aSvmxw7jLFSd4+WYt4JhH1EQqkvr9nrgTPlDw7UxWY/zeKwE/eT
MICUT5AS+63TV+u9OOAwNkpWZ+HgtLCAWVAcdOnuY5y7Te0Pd5GUBq1mH5r2tfcXr+DFotMlUb06
3yPboDvxm/W9YQdpJMk7xJJAKMb8DeJA0UtyMp9BYIi9ENmEWtuk2kF2KkkkqFLAViupeaNW3xQz
dinBzo7coM52TbJmbH0y2uKaxYvIkoWIA/0PLQGkSShhwsWj+9jY9ksIC8faZUaaHBLWfI9QDlm1
iSB0wZvaaGj0bEyfhwtQD1bqkAvUBGAl/ykPGvgl5JMXI/8k/BE07d2RmOzdhBRpWQwcb/P2yUWt
Vms+/vwul3vY1pgLGWTIelN2sD3U+ZVzw/jQTr3mHeWqaHxd6n35c61DzpU0zjkMFrqQOCNnsuVe
k/G+WmuNYC+dYpzagtWMn2ZA1DfH5tjtFUiWuIdiL5yvAyzUip2JDP1ZMuzhmbXgtMYDlkNndIQZ
3ED7jKEdM9MRyobeU4THH+FLr50pTXlKOhwIzoLN27p0Pl3VgHONCnW/HVhfo14icEDsd86eF/bt
72xLi4ykj2Rud78orPpVgvOr08nvdcuPqw3atUi9O3NnYN4z7E2vqk7uDLTeTulhEEjg8h+T07V9
a7RFa7yTAnerbWaJhfxqn87fZ1eG+5mpu14cGHtDZ8ZXG0+UOrroxBQD/7anym2nmPQhzrdInK6Y
0TOEZl+ECzdRobureFqTZmpMNaDDaRQMhXV4MpLbyka5QsGfV/I3ORqiCK24RdBmTjo7vn/5EAKd
FlDOOSNiH7aNbKjIx8lcaAHQWLe8GssmEpC5bi2Uu0/HgVU3TpnrMyE8icou5GRCeEqcQG9GN99+
zyFvFgpE7iD2WsY/RvJwToOlDzu3sM9fFiGe3OHCS2KF08UgqCjcvyCKfOpvxahFn3VY8oXKcEMD
/9AbiElpQNeTphR+DpQQbdljldbvYAC9UqZND/XfF1ggtC7L3woU508Wxjk1TdNBGEmPJ2xYNnkI
lTrdF6bXI7MSeOhnp7EHVTt8RDktTlLjjQgaFCcxWzUhPLXiLQSfMD7xD0yDo5T69IdsDW5CuirN
fDlViNRvQ/IS8xk92r7OILzcJlU1NFxJ28+RYitQPtcYilOI3kX5eMsI0bFXHRRi8BHrMTpVUx0D
PRzlC8lDCUgAgxEsoV5qhKUxA6jxsiRVG+YDcLDPrt51gD8Jx9eYuhOlxUi2gmJn8l2as+1M2AGF
vFBZNoPHRVE3jB6LnNykjHX+rBPtKAfhGqBEQ6jRDhRI9cMbXv8FiHs7KbnY+KX6wbkJ9bbVc/eS
Mb0UmOXOWBzNYsE/6lPCLBrsUZ2c5CNdSo5nezQXwl3JLRx2lCslkZ/VhZnyStoGCrXXH4wP4lFY
8fGR6p4HEFdR4nu4b2eQMLISyxogFkLCx8yik+oNhOKa4O8CLzVwOs5yX00l6XYWlWhRUJUeMGHz
vcUIyRYKh/m6N0DhFjaBT30fxfplX1irZQc0qy3HQ1dbyEUuRUA31ql29U6oSwZtmcPRXoc7XxSq
54KqSsO7rupckNOGMvhlVcnzj0RTuwoKDUeas6MZ0ssMGcSSLz+TZPUmDC0snGvfNvyQPwzKzuvX
tUHc5D10GpeMs6QMNBQiFX/G/B+iGZQ5kZaZjDTcrFzLfYKpJiMkccYu/QCH1hqZ15aOaZ6GLucK
6shth3lKsZatINENWBGUwTtPMELXxtInmJee8knLuNhUDYBZ323ANE7yTdDrBIfuuRHlpVWq7m4G
XU4cEh7mEDyoqA+sljPr9wYvqaVXL/m+f8rWioLtFnInwliMmixAIMlWIadJSarU/adSl/Jvs8TY
SEMRbBJs5oj4UflY3xOgRiwxGDCqylgBUYEDSfq8ghfz/7vSJvij3fPV/lK8EjQBbeqYf5NJ9gHs
J0DRa/sAMz5wDnyyl0tkuIbxsnvb8sw79cd5cGmDysGJSYXx89axKRZJ9kDW7OphKdD3bEV7HePz
63NT97YHhSAolYJCIDCuM1k83kyVlecXXuZAA+ECIIm6cQvozE6edxTaLCZv4/oDnoMfveqlWtLO
j/yMWE5ZZ/d2QPeMWQ23jkjfI/1rT2d++agWHogFRcj4ARoDffL/3TFFkEIuSRUj/wRNW9fKZpfm
xBv9bOQHq7jJ9PVl5Yvh7uKTlR2OrJBRbzVBc/pc3n4/3C0OsCOtRLBhJ2eOlKrkOK6bs5mk5tTX
3DlmKAvirdeDjZet64lDbl0NwiS6W/gov9LjgOgI4SpOod4y84divNPegNI84TZWDA9n80qJWcqr
FGvWpOdgz6R/XLY0sbxckkcNutpUaoadUMWL7fArQIJ+QTVuoBpKzs1iXsu4I6CWEFdZFxOQ/bfe
Jjnp6QfNn7oPH043FYBgE/EMPqPMrm6sWjmD9zEvJ0MPmi/ZXqBwMXE31K6SyRA8WfKxx3uW/0Io
bfLoIzRuBMmwdm2YiZFiBXpV0hr18SCo3TfpwpSIJ+eZZHO43Y+jbmSxAdJjIQPEIWfN/9KAUbZu
jtCn/fNcnRQNGlOw4ufGFYvQIsdljv7hvMijPzJL+mtRlwBC77jXhDMQEFVfPkmgjRXyl04Ah+Xa
WuPQqZRiMg2wFukElyMg5NrSx+7Ri6I/MQUfvsRt6QmQwZ1tukt9+Yo21XsnoO0pBhbY9/TCrdlZ
JqO6YdZYOJRXY7mm6TdmZOhwFt3o6bucAGxg9fWJu2ul8aBk1cvx+yNFUqBgs5bt4ERjDRYE9H+V
ahZtm40VKTNNuGecxEmKd/dJ+9M7k2Tk/pS31gYQClUv0TOcvd4KYRJS4PS+yyul58+1Xw/VCcGs
scR8NRwc2Gwp0F4OPYYT4/cosqfg2PhdEc27zdnQM3b9XhlF/v8eHyfJyQT685iLb54ST39msiT+
zcZFQlmTtotlgZUvhs9BE110Wfl0d1w2giB/+U7N2Vt/mfKbTlvIfyrd1J5R1wcJ4gmMXyaTA3tm
TGibvbvb7zquQcTkMOvsa/Plw/pVNFvZl0aouEMBwr2bpBtJmaZUrWhQME6E0kPZlAZUCTkv44Qh
Cjrgv+qoSOChSKJdo62Mt7+aV4ZbtG7t0sTL3iz9oIRfR0wT4xuS7/w10FUk5nbMZ9Ons1X13JEd
EUXDlw3hT8HvBEbKi2Sp9knHU5yobphYitpQlrq6lq+rl2jr88hhRmZ1G98uikbYwhwyY3M+AU/1
B1IHNUdYoD2t8wtIcj82ubgbFV+LfUxEN1OoQI3snI07b5QuubuwzPRYAULBxq6SHPxgvtq4jAJg
ChP8le3pRNxerEYs8LPvA3U3tNTVu8YhcBvkiV/xlsAgpDmxB1sgLuG/axV68yIYQx37XbAZC1j5
UeH2SpLIQ14BCtxydaTkXxCDzbGsYClYHjCqUiVu/HUvEXeanvZpqvSE75SmxydBVGmJBBotpG0p
PHcwQxOVscw2Tsy5u7+NqGzrcKeFNfwhpps48wKY4zalQLmBotTKkoczQw3wC+j0sqD5liILivrI
P3ri9mUqxWdX233DCFcF9DRsVPlmKd69f1VrhX4ttwEGinGegegRUIK8Ofz/fRPv33AnK1/QBOY/
y0NCdfSsFZ3p8gQkSgvuAEJdNSAZiZLtcrreSi/QZl/8BLbuPe0AEAur2/mUCd4FmKQVcYVhf9aC
UBdx0Od9FUvMelmI945CLR7NAYbo3QPPI/i8rWooNjaSw7ioyj8kn5LzSxfa2fAivyOq8/KcdnOs
LlK9/NNt1eQtQhNUGYixUtnmEWe+5tz7V3tkRrHkiYO0KhBb+Aam8Nr806i2Qj4yFn9Pdh0zWk8I
e8Py0ALiVbVMn0Mz0jv8MUBcoM6Cq82FFrdwy6l3ahcD5xzEFG+xGA/K5bfndGAO2J3qgHViKREC
gI9BkoZVJs3ZIk2byc7S7/+50ASyiz2AHqaQmpZGcmsGPMYR8ZDM4wPYsIS0DTCiFcfqtLo9+fpm
YD4i0wGC+pDX8SPydD8GGYyWwhXdWuPiOvgr++SOgzIhM3UCrMS1ZzQSMAYMu5pK2XlKsQKYI3tC
9ZmxoIuP0Pu6g9MAJ+QKWsOxbGCYS6QFXi3O+FMbkD2RJMchbAEHxdNyRWewP0U1HzP586zifL2c
EsTNDQnmepYRQrRgtZULdrr3hC5NwFFjYM8vfpDxQ9Mvo1bo5/qBjZ7+U04EzgKH1lgtDLqXGq4N
2oP74GjiGNc3pIieN02D1x9+3ge06wanGaGrGATVfNaIxmUuIXy6LgEcNdD9qrRKRSb5yFJW+r8e
Dbtx+5VVPfCulwIGxN7o3aED7d7pPnDBYR5U1fjyLIaro6Ff+ZNf2WkmU1RAfVtUKAyM3C3QoW7x
bJst/wZmtXDaR1GdTAiI3gYCT8jfHkU1r7AWMuuZ4LKQrRlcGs8xPvR6Dr7ezLdzKvqyjH4acb/x
E2nsV0Fs1pc2wp8HHKTwMMNXHGAMViO72fDbjR6oK6ixYttNqmSL3EoPoMoTVFLh5RVMyTxxzxFd
lSZHuNpmXa9s7QD4p+5ci7V+VppHch1x7QgzI1hi1dGcJH4DlFunelWFi63D9ndHKbTcMII3c52/
QQbDP9WodD7eRj70vkveb8uVrqljWz/BhfWkFds5SQbIc4rNkRd8+vkv/Kj8MsRVlcQh4LrICoVI
N8MJfcmri5GicHV5FTa2SiOTsVv7Mv3X1OeWt3RYLR/RSpO6GJ/cqQIrI61937y0QWuJm/fPGoHx
KjIFvgYi29g4pG7eC2xuEl6Wz41fEyQsGjbtHAHTd/VVGG9drCRNjOIsm1tKmWS0aR44QKyxA5QA
tsAhV9uJ/3Bvf9iN/6YhNSwoYMcOt30NgIxV3sWL7cTzDF+tUa3BE7KmYw3Sy/+7GOXtY/v1hG+U
XKCFflAzKunSzVngRh7qSt9HFLRzqEkbd7O4ntRMgaRuc+7JVRuKtEy674uATeIQUAEHNilMOIO/
fxdO5ypsq6v51r0ZlVgoMCmqzjx/jrFm1k/D/ovIho+qLd7Mo7Jlcb7YuZraOjXH947X9OMg/AM2
TC2saXkrm+GwSBIF+zoZbPFeSSWnXprx008Uv3CenebfPDzlo91/Neb2IsMquhADNzWenlK1CZod
PneUuLWtzuNx07V8RFq5VDRq+7z+VDwBixelySi5FoSk/gHds6HWrTNFbXkz+ynUIih/wuDmL2GD
pVFmdv3hwwFKfnO5ad9mg6Uz4DTmV9lLVFXkg//iorucUarALqfG7lW64FWXVPcVMzQvi8/g+N6a
ow42L0Cm7Cd0Sck2Mt1OIejQdIVVTDamhRNrXjKJtS84s467m5MnqbC7MLeA/LuA7tWjzKw0qGzi
31sS/W6tqKgK1drK2nH6r/2i39s3pyB3L0uAGl31qsL3+9Ly7i2vMNh5H0dQmRZaj9azH324W838
VmtSiuTcsXszADIKmycVWuiIF7KEEg6wPk9hDeYacgQuKbmNBVMEObG/slAQrXBA4VPY6cZEMBE0
PCuj4EDWiVULLFxYVAcY2tKZHQqP1eBv/ByG3auK4A5llFdgEATHbnP0zRfzxk3PpaGzm7dlgHUE
LEAqhXV7CCU5BmogQZQHSJrJw6CJ1qflj5gfAvY0KDqOW8n0wq3RC0iegZ4ZVjPt7OimiJo9tUYz
zaLZsZVjkybi8qr/VH54+/In4Z79oKnMnWgMYQFi+FkoDaqIwQUOm+6/M5qnGrGZBnocuBKzhjKT
ig6tm8u74zSUiiyE2yraspGjHmjvkYUUuerid/MX6Dv7oHLX1V9+MhWXgjs5XbfoIzkwuBlUDTyq
PGKruoJlHceTQXuxmt5laW1XrlYIf+TH0ApEcu2gVH8tJy8nnRONNHPyZKvX+0wq48IIYC96cTJz
jj8ahg+CNGFWeE3a5ZWfkRjfaeMXRjvtYqEDmcyWp0IQdfrf5K8z5aC1qAFdtluz8R+WN+LfYAqk
IjKXwKvccJsRZQvug+8N9nBnsWWJjmL96Z9qQsCtrNP8l5v1O0VWyF8FKuHJezJL9LrpFFebEBUw
9FK8kNwm7Fw3c2LFBEhL26p2F0FGAs/LfYp2RqPcaVzzxEmfMeP78LreWnbhGjg1rEgD13ZdivXV
5qPX965S7nwNc4z7G3oZweh73uX/pr9t0xRVD11s24/rO7kk2gvVwHZHFtrtNqJhxKFQtCK0nFC+
ShTtZWpUwW/q8bXS0oPZOBdjAha6Jhtz/I89GI+otBaU0DftcqlT4Nd0zkq6Vdfo3jjIayG9me1e
OUXJ6GUEx2J2ats30Sprn0et+HQmZyq5mQ9TCeptweGAF4AE58So+PMN4QKRyVHyP8uef+ktt1mO
Fxu8/Nvi5yhbz+wpa7ygxn/2YJSF/tSKXfZY6M+mjIIJpFiVAxNjBr1tJ4U2FfQmp4mtyRqnqP9B
94xF8EH9QbLW2wcFlCzR139i7hVy2Oh8wXT9/g5PyAQNFHQmErolwk+02VnITdJ1EiqFjGmfBPFI
dCl2sTO2cKrOi/BLw8QmHTFhtNGNuupLnsxn/LdupBbCoZE9dP/tabIYUYvNgk278WjzV8FnRCRC
nOPucnqx0hT4+jvEr1vAP4nL1MHHaJBAhVOdFDgasPuMFZCqk7XmICCUjQk3k+dWiI33AFp8J/wN
97oridypVw45JyrYHhj3imfq4/ZL1A7kq6bQirxYepC1KyQjiU9Lqb0dAf8P6nEehpfBx5sldwML
ZjKNdUKkfH7B0sMFaacEx5P9kyeCYMCnIUozlgQueBh1lXf/A2ORjg/NwsXSQM5MwE1oJpZSOkUk
9fIO/g2VIJUzxcUP+N12o9ncMBQ0MtKuqLcG9rXk90kC7WSJzRg0v4UcqM/lF495dF8s0f7I8HTm
Z4bZpNiVD0Pj6eIx9Pn+mineydG6jhKgaDuuHo6TvKPbFFE5KtyYRiwfVlfJ5bgzAv9C2dJmpuij
BnOXT+9G4Ty3j3wNa+bfb/fwZgkwEyBahPu3SIR8Y7wDKgN+3pXZt5Sygw5x31WUoHmDvt6YHsjl
Sr7rq8OF2TTTHBmzC/vw5EOcszK/Mz/9FONq3yQZcv8nYLbCl9abZC4zH7DjDWa0fXfFMZ7nm2p4
aRXUpvFLggBRlV6nVoXhpD35SN/hfP6sG6gezuSzVbHYggg0eM9dkgXA9u9qm5MYv8a88alSN9+B
Oniz0k6cAUIVJRr7Fg+agtPeH5Qdsqrn2hecix9hSwlqfyFqL3A79DzKJ2nQtm70vh5k+YDYwy5i
ZS1J8z582vNJzPneg0gd8OOXa9SD648igP7JX8Liwk0Sjsw7sHhoEV4p623JsZFjt3LiPhrqdbCN
phs46PlB7Xm9XG3VGUEbNZLs1lSR4O9YitwQ8aPN3QJtnQOLxprh8tnbVL79b0vefBKNsLAjrnl9
u3V+Vus02NO3p3FQngIuZl9jqGnrw56rpBlUc24u9ppKdNGk6MD1fFMBb21WfpgOe4b2bdJlUqRY
ao4jF4qfaseibkhRaEwMr+V4Jdng5v9rJmA5w7zrJukvprTP5fZRcn2WVsCRMJ/gDR8z4sDcZ6eT
i9UQ8aujLiMAfAMUG2Gs7H9GMLVdeSADJebIJCG2VWrjwEZbQEUaQt8PRt+u9laVdiapllnHeOvY
WDLtB/LGY8j9NQ86FgItvTgPpq5j1ozDej2oXhf5GwHLLJnE+GVksPp4a/9sBfOKZxOl6bAMP7Sm
cxD4gSzQzHeB/9ofFpgHMkGH/CkwKvTz9naGpktfMMm/UWFkbD5boaf3OnGQFsG0ozY+wztkox39
x4FVgfQ5wHu8nhTdKc92+frFPEmnSCvHoVtBtkXoPM4avsx4WLflfoVyVJOTzDySw7jkztww+13R
dzgnmHYuuziDY6adVidGP+T19+iIk25aOc04cCRW9uuhc9+fJWnG8WdQaQoxAJwNrcAuZ1FSf4XM
jtr6RBVXqCG3ig62zf/aHCAXQt306S9iN/hUiVYjyxLLgjVKy2xuxQygKzCktFgDjZ9jj5KL84PW
uqo9IMOED6lt6msIbY+EmOFI4G52qY+hZOWYgY8Q7O+XBHArhGOcwdpG5OGldbZQ2mQvFlGOePi6
VLGrVZRdsph4dIN98Ar+mbNZiqu5MeagecoVcRM75KfG+/A3mDuJR18vM/wH+NxXBmcVONlSoYr0
GNYQC75hEVCLmwjMOJLfA/yd7+tlGc9zMX94q2xmQKY3umWHiQ5UGlTcAzRMAlJSJIi2ieb8mBG0
DlNi1e4McERxLzuqBN4/hPZCVt2Ftv8uFDiM10ZPD4wVVpxkSdqSPOxXlWLVLS+zbczNEPNSL1bK
t1WHJR2RLReC9T5fFT9n4JjNnYppuJRZM1frgtAxdsPYDHEIRTWXcfKqDQV9unOnW8C7t8KoGtCu
h2vZv+PgNofRJcOdJwVkmHnGD8k3kxtYhCBXD93k5FugZS2MCs7eyPkvkup4/2GXYZcWNQSJBNhr
ZbwUTXNiVR7JtThIxbVnvBFe7GOi8umw9IblUtyzGRd1gGXFztXW+UauHQj8EIGsgybGd0gKA9ts
KAMBuviNU8TguOx5jK65JGEOHK0wOUuBtltm5WeDRxFeOcw3MltolcXYd8hQwShEmIzLZJJrbFgw
AhKnnPTQ78BDicOB8dJM682i7lnWMZAjBQLBlGI6PlcmNKrz5s4sdZQh0W2BhmheMMiAj3jFNFBX
salVRNCvezaMg0P9eXyUqwemY/U6FPEN+Y3So+aTRKd1uY/vBgM1HEfX4r4hWQREA/3I0b9TcLK6
1LY3+Ze45WSzODoZBeVjgsMEUXSSEhIhDX1lmYOgT0o+oZvOk0K4b5aHKA0IZeoW5niqqO4Fo0YF
8TNGVSPr9DKDV4yYXH9SAmPuvzfJfbxMOF8+HdPsK6GFd6KLAkacqIbyWDJvaJftOBBKYYIaLHZz
bVG1sJBDVFcughTuAdUVTUSyx59nmMzAz0I3xw4LqoNjYIujUOhaaN0F24A0HtlLHUoe/61gYYI3
YJeI8wRKB1IZ5T/V0dzeyBfJRYH1ykUr4g2yDw+4MwrZrktPbfjdPgiHSIkieJpjNCKDcBMEpJ4q
g3dsy5FudyQMlrzXXHBVl4NBnrUJmAPB7eZh1/AKTysQhPyQs2/ptbaO7BeICI6LwFqvkyHPfnN1
EUosovN0BdmtL5UV/5yJBhrMvrj5ZoJmx9xRHgezEhe4ZZiDGQYTznW3/hxWIgGkYTf00+2aze3s
GCWvCpARNawKUepdiW99vxZL3Hc3A3OcKpRGqvSEevV4o9eqXQ+MiwIsTPXykgIpzB3mvbl5024o
yMQeN98uFH6eFQ4auyhIdQ4hfVCHuxTC081DUqr93HQBc0KC+2LoYKtolgAyAMGP9uoAY/jW98lv
ACkdMqbCkiEorMPA2ORI2zvhw1PQEynIucBDfFMioRYg+H4G6JL6PPAftlw7Wbwjd2409UgdPTzY
aWdGtDXQuJ43GzPnsQ9AhFsy1ZB4LGwc69NGOjs11LZbQ2UJFhOHllPr7RRVW0cxFoPnp/urT51p
0yomAWf4me7uRulmTro5BFYhhCdXZe/jdX9NJ+VY0Sl8/q5kUoXzNiVLpAOBqDsyD+Cavwane3QI
gNN+bWNmXa3hBFHY8Jw6ljJD74ENQXtl8dqhNbTtXkd1O56gfzcn/HkBStQR7YachY2cJfA4uzvu
qgz7Jr2Q4N5o5ZV5LodRUpz6Vw3jEbTLEgqDK/2lIjd3FcC5WbMplrwJTYGyqz+vBG31uDjn3arR
EnrpSr13bo6lfAYADuetB3twhDOZeKzqAFHV8V+jD1q6HVksLYhQFjg6HCQqMGEWjwxsXWv4u65v
7w+TLOdXRAtHg8LFrvlirnKD1KOnWlkSBNAMmcnTZ90vN8CMD7azljf0dMsy6Q1mTljyipI3Bp5X
Rx0JYwTk1+IWFdNQUIheVN4nIh4L7kAqj8KTxulTxhKTiwgsXtVknfeVsJIeK/SGiT7JkVpbZLv9
I3P0RqY9J4uK2Jxr7EWcXzOMGL2Io3xfgHFV0OuB603KIRdpMDltyd7yzoxWM7lfn05qmg3FKk7i
VdCj54Ak2fPdceNyb+k0+SFdShcrTq5NjwsEhEtABIynyTaHKNtoph/3hmc0P4xCGc5ICVWascGJ
nQVprD2ogvdn0a7Brc/5DzVUmqYoVeaQ3V7ikLu6qtaUCDkqG3+m2DBERoXt7oVqSJk0J42Nd65H
RA61Pz9OGaSFMSjz6rfQb96VtfZ1h4Lu0BoSctJUxaCvhXK5smuob8VQI7jDOZHG1ccNhT/Aytps
JebPjgwNpu9WqgUFNRqhLpY/c69ENHbrsQTd4+OiRF1LjoM8KPWE6UeIPSdcgKqGpmtadDL17KaZ
0BQMyf4BIC9FgG61ZXZ7UjgyZvk8ab2D4jAuU4v6CCTid9LDEV8oqkz7XR69WxdwMZRmOYCPLfn+
nFRUFZVj0fKlP1iLfQHTJPhkmRlvbYlVrBE4Ff9JHsXuJ0TUObitnMAziXhcGPtQFx66iCXnIhl7
+mffkrUoK8HSv/7pD42pAqtMdmjPE0NltINddGltesmGAldyflDLhnbasyJsQGe1fCZ0LwAfH0Rz
YLJEH1LXffpt46HNqHejTIvX5Lbuas6b+wGedsGnqIns1ZaOLPgIEqb7VAlbEeV3EDXWcpGm0Dhv
OAneMwMz6ClcfySn6UWmuH6K/Hu5ivVudKjISuEK8lKynQTCltG1tUC4wfn+IdKXGBo9xB5/F3mQ
EFwbmuYD5/G1X0o3AGu4bAKbRw1YNUAQk/a4O+AchMTp+XYzKe2igsuUdOZh0SzV65iydKULGhoD
1Xu9RSXrmKmII5g8m1OZ3EdwzZk6Mb3sTYTZjCoHAfiokZQI0eQUoRfEpMvwAixeBWKKbeVbIC6J
GGuHFrmwIouQJzgPRCqcyZsnq45v2520pXBV5WtN0pZOi/tlYzk2dompJH7gkeB6supEVT7GxE5Q
bbFkTaVUFX2qONfJkOXAUKblss+XLLIqxE/mbKkS03vLjbQPqAQD8QmJghf4OUlPzt2WriRWuBuv
aaBhqqndOu2K1v3H2Na5xsIQfgBax+0iC3KXHe4JRjg++M/mCTQ3KtXw/gmDi57rSeRa6TIf65j5
zQqE+gb3hhCDB5ChgxIjAfjZ4OERQt0lCT0hgZ+vN3b7cRRcQms+xl11q4Zbh6/ujuuuDaR89x/Q
G9tdNzhl52OhwOp71ZQ2ONCCBU2wSdLkZJ1ZFECJq8ov8kvBMlRosuZGjlCRqcOZs6ErinpLLrsO
jvgjvAuPx+ryv3fcpIIGQ1fxngwDXDJeOoZAtbwsGkdP158rAOM8ch3jCygzsrXR2UTFV7tq4S0t
bqHWfFs9sIS3vdyX0URfMbpM+ZYjjUsaEkYDfw512JA9xZ/4cgqejdXOWuUSgUeTK63J4wW9Biyv
QQrMxK++9DV5LodgSjAC6RpwKBsk6DL1znM92vRJOYO9GMVLzA/Gid5pdHtrCv+dxSiYk9tz8Fxt
Z2GJ2YrfnmZH/VnOi0JfJGgeWKUTTAdTg97fAvJde1xKgBldGFFlbdFpE02shjS5uPtQGOmT+N93
e4tZDZJq8kaqjbE8VVyfFe5b4dvC5mlB4uQTG2o51qmRA2kCiF+ODiLRgBeCvoZETvGllm8cGosF
bNpVkbJeAV4HKybhJISqFnG7aMkYlkreeXaeXIpkNo9x7wfuFuWwAGvGG7HNTEoAAT3QSqJdbpY/
F+C0KcsOui1l2n+kGTGBLvoWBDaeOP/0AgxDRfutw+9neiDc1lji2NYzV1YQXt6JHPiUdT02VJdd
jnDcPDrcMHXIzulwSDAwYf8lGGmlAil/xMx2S16OP95nsCQKMKWQ66hLyGh2I5U2rumocsZSzm2X
tMei2GYfjPRNX5MSi37gGVB4eUamAo+522oWVKtCDGbThJAs851ajI2up8Qsg6ZyLdh5kxZOP6cI
6UEEGZ2f8xliKP0EXwyolp8qBGDe0pAspUUYNOebonI1wVfxzw/Bi5590vxBdlh44h8eV8PgEocD
zzm0w6Utjq8CH9HPguAehzGbzn1PiC5bwWs8f99Fz9ZQtlUorLs/r/c/7QeSu9IxsW7lWFkIq1XP
UEbYdjw2G5n1NzWZ6pLY5yqJzxiMoEnKXCh1IwltrAWzHxe78oKuiXCmudLZXOa4u/j0ls+i05Eo
9C0SeJj020OF7Wg6VWKORYPxvaa70FBYdwwNDjvZ+rSj0uV9TyitbH7Cy2JBjVDDtOjeQG5/em4y
+r/w9lC6DoRzwRneZBkWhNS9uBpc6WaZBxewZDj4uS3PPDEglbTd6yZDq2dDQ1sB33L8PkX5doV9
rH7U7o/crOX1vkUHm0/Y+XKFVI6fgdLMbWIvuQ9wE1L8sgqhggJpm5kSsTj4ZCChUFGFjfkjjshL
tcSfzcWM79hpN1j5OAurE5SxSA5mGtDWT8KtB0zb8sUVJKPWHD3pwoC5SISEtCPyZBXzyve3Fba4
+hn2SV4kkePNYkJNCw91dCrrr5Ny3LO/JmKHWSGCUEiHbsuawPvlJ9NWXttA7y9O70LLGQv8f09v
fE03Y48kc5tNqGDwNTXPAxJ49oby2K360OBXrGWtBzjcaupZy1Ehbd4/DXGbw/F3OJu2JrTbbuG/
ybeFfZ8H1TneWl9CywivD1oHBtZXXnoj3FojjWaAoohylpJJINuBLfT0yirTJHypJNV8JSAoCLAQ
XVtUjVufcT+luG6hl6qZzjqjXctE3Tk7aF3/P8mecLVx+Q3VzqKSiHgFg4xxOMBktYZwIJXM5cw9
9OAVjZaU3hC7ty4MR8HELLYyI5JBB/pWrKBZNEDnLNUeL/2y7yzX4XUuAXRTewhliz3THgcEYjQ7
XEs5dZ2ZASD13vrYQk1z2Y5wmhDzzi3W5wciayhtezDfwYYpGhj/iahKCw9G/bFY30esnKt6NjjX
ONdJpwi1ZQKoAFdZur/STy6ZTUsdbZ69S97FmSstdxIztRJi1UzD4Ml7BwQxlHzj1o2x5UguIw/h
VifLHbjPFhmxzvie7cqxooBc/X+8IeESr7eYUeB5/+qBpfU75GAUGT9apL7Nq2gpbykff6QndCk6
rtioJ88WfSjRI8cfG9t6Dg2tR5sk4R8KeUA8ELZG0khHLvklpMOH0QWYMe0ctO0T3QNSnIrrltge
vV3/6iAHMFT9RIiwY3j0woUYgE7sHVpKSE56CsxYyl6/lQHXtpDYFT1UFIoDZl/spvHClCbI/ZXc
c/9hgfCt5XBHPN4zUtOdVt5rfx+8eiSNL8kgErCRRn1N5oj1CKlxJ3DPFvnugj95qDvo6lb68506
F9dXEmicvRqV8SY4C2UKaQ/c++KilBAANOeW6DreyGsPur1EYeXMr/GooI1ENyp5kVge8oGguvFd
omgM0gIIWmpgGoDl8oEcd7Kqxh4Dcp7ilkrJ6tWrW7bVyIZYV01d/jKYa1RDHUt9MIhSaSDn4Wjz
xA7cCiLAySWq3hhcOZUJYHIVoo1pWxgRb0uez9mJy7PGvjK/zc+ntN9JlRYFOWcOSnjsl2RQvwat
hN3Kc7NRVnqk/SIPPEkcg7Qhy/l8k2X3jRTi1WvlTNstsqqZlFmfmIz/xc3Nd+/LgNtbcNFWTaFi
cQpawvWWSKBKqQK9a/OX66kQgZOfbIwFwIwXGIPbMvUyJZSK/3VyC2vW3MBQAJ5J0CXYc2e1hS3d
AnOI65t0tNKEDqtA+R8ZJRCaD5g+AucNROzaMQ4RAmkyWb+fizKvvbaDmQbUBnlw1/tux1j5dCEv
qg+ln5LVeiICJefkOqrm48dNWLubr89T7Cvsd/WYctItCs20BhG6oOwx6dDvGxdJpS2utPhFKLiJ
0XDHw+3B22fmuGIh+YxpJWCP0lnvjPg+vLyDTZXBKWn5L3J+bE2fOzRX3ZOPiCFtpMhBeEnaqMLd
8M2Tqj6RZzAxUapgpMiEOYCerxK4VgW+tjslK35OYuivSJezvaEuUlIktIT9uZ2baAdcw2kJwNWH
ktCRwSFM/sS1zNPPkviDqkkqrm8VDjBUWoOClk2TK9BSoUOA1mfl2qoKYy9VzyjsfajVLBc7HrAf
K/XPZpBGTSQhp8NKErg2UGtSZyBH9N26dlcDu/RY3N9jDnTCXXFtggjSmD444CgqIS/SbldcR2qZ
zbluqZUIYjGrcxsUCRpKesE24IPsHVr4A6IaYTMe04OGdMVliuk1ixW8f2g+9MBYySMAbGToBdXy
Ly7yyyvCwTx1qqqgp6v2u4R7yvTR5NHOeUBY73KMhKHRPHKBtbxnWDZHr9pcjmh9W18VbXp47nvG
Ho6Yu8ksMjHnLI9JuA/wbKJEkHc9EvIY6S9PK2b6Qr0mR65rMeGP1GYmD4gcDPz13g7TaunxTZfd
nXYw8k2yDi60czs9xflbQSOOpOBuQznWrzZxisBqK77QkG4n3afPsDfksN17oBrjZKzxh7OAAQqE
opi1Gm5lJkrSP0BAWyUs3gWEext/f/8HI5q4ycbBb2iNs2tRhqLClxIFSpAmfx5RZIcmS4isbUQP
0sSapXSWbg+8ohVycBMSfmgquxgGu+VsxfuBFf7CQmJv2hcXLX56ct5Oatw5YSSjSPzB7omJuwgy
wFVfV/0mfKpIRhpYnMZvm7/5aEQ8ahVZF6TRKqgy4oksyoElK24LuZYsivZ38uzrkS+lSVFhs+vR
xuvt7VlJ6Hn7UkxFOMY1r2lzQE+UQ6a0b1ODkSA3xjiFBBq0ZJZfE6zN5URyrpB4F5psZh7j0hDv
aKtO/mkGxD52A51sBFqxxQ/c37r85tIOngWAWS/jAcFd/u1FFjxIIMDGVCu0AZNQRyD+e37GI8df
DMbM/PBsrK6EGRSXsOrDNwxtScZ5UbUH98s734T35WXLTE7onDjrNGZd5N12Al3vY2OjtNZYyV6K
JCdNofyzCOYiv+rc4YEQ2VeOCfLYWcfQPBxgu94O5sMtjap9lj3ulP0WwbEdzEBShf8YOc+7+yIp
luHXhCEFShBiKldYSbg8FRXeclv3OixQ/NEPByu0Q43XLFvvY5L5OlXQno9niwG0bWN4tsX4Jbt8
7MV8WzQZF1foX1uhGEoHNENQGQYfs3iAQugh0zZHbVu/2qtUSNwGtg2jjo6EfSRYaaOZ7iVs+78o
b5kAZDddzYO6p9xU36xKMbAYFB4/a+VdjZc0/8H47plTXRee9lqS+58hjQJ4ljgqfz/DZ7eNp6SI
VbRuzJzFjvwV7/UH4oJae3+hhlMyr+J7O68Qu98DZbTNr6AVPM6+BAGYadd0UkxgN7Fu63NiEdGc
lBrMb0aV1Qe4VphC3nAqjSgyPZ25duVE0b5mPFsLd+HBbU4bovYzZR7ejGa5BU9AyzG+3D7l6km0
EEH27XNfbBzeM/TR8O/LVMt13Jg0tagsdi2eb0gmVXIxHtMQ4V3oGF+NW/nPXvoXHmhvWgCEjnBx
WZ8iUTdDOQj+KPNGrDccV70wuQOUmoF0ffvQKajrgjjaobU66cAo0OHt1IF7qRIxcZBIR0Yxxcqi
xcMW4YN/Fes3dX0QxDfgw13OXsyD2NjypxTljMCkJUZ7Oue1HE6VpZRX00F1+9iUMC/ykE9WyKdl
ChOxEzXN7SjHyxHsPWm2pmR68AoGyjjWlU2C5QBDStv5sygbpnSPOwGwK/Ke33+xh/05w+GZzIfi
atDYO5ASJvl+LzogUWJZztgWVV0QeZtp61buQ+1rsFQYqEfWmrj6R/JVcWLV7tJh8x1hD6D9ySUu
UZcks8x4JOLiHX/xZSY6+hhEH6pN7Ous9pGCDXvYkN2yKm9IjNjdRE6opcZCsW1DbOln4x+Km1Kj
aKngrCK3SOosIWXaK8fYlvQwkipqvz65dj5Zp97LuVdfMfcDs11NOhpAnX8PbiqTh30QvCtCkkci
31h5urdub1tzIK+YnHGkgmkwBgMJynBCErmYxnwu0hFZg3Bx3kPHUH47KsyGkERTJmfaGroW7NsA
8urw9iAE9Pu01xurtenlMcVja1dsqCauiZjftdc2hSuUebXMc3iFp+bvGydJco3kqt9B/ld4eqTF
C0vtXG/WWsFm6VpJOwYacFtRD9aXK72uRi+ZPlmsqKy0NlNqlE87/+GUk8LGUtOe4EmhO7T83P5F
NrHyWxwVO4p5QtFght63rzOjz6zFmZmJ9q5ZYgetDpO5Sw0ikF+mZmIP1/7oy4LDUPcR8uL2G8gx
s+Q8lXdUGQM70m76//lrU8zCnEKabtVl191cXACeLo5R/XaZ/+5K3GcMIuecD8fue4ThTEcaTq/Z
TmsS2BoED4wDhfbyMKxoNBoE7YROByfGMyTz9lAf2Ax58/s5ew7X1GAcTgBD3ZA5EqMEP3x7U9mm
gmiAc7cZZHxRitqKnords7uSIZHDInzKVLJ9opcyHgplZI8mrIWhzCdtdcXNNooKv2FfxnqqER/B
rlMz2joqcl0Cri2I0MLnTLOO9faVEfzYTz4i5qsC8XvzzZzR3uA4RV7ItbsR2MRdg9qcq5NC33UI
Z4jbZtK9nEI8CescezgJHV4ui7nwa0jGFIxhqtJ9cXgCA7Ie0+LguCyVhpzJC8MaXiB3qZ/NP4UM
md60Q2P7wz+Eo09SMsC3mYyoeVDF3FuqOGby72265LqmlET5IU57NVOqDbIIQjtyyt2gyIwPnw2G
G1UCd/fVmTUAnWITEfTcFuLU1RwxACKIqv2r+aoZLbGZpHRHgPAzAOS0jYu6uasCY21f3r8DLsbk
UoylCEwj2xK6uWiXkZBYBHPjRxaogu/Koaftk7+AaimeKCzdMzkCHRKZu2AqUE53vp6YnS8eXCuQ
L2f/ApnVg4vGK1mji/cXY/gpMZezp4Iztg5qDysnRega3c8RDNDNYVqZIoK0zpNU6eM6jCOrRIXS
Un0aMOqIAAuf76xph8EE4YgtP3an+yf5gonqODvHvwM3sVvJCg+9TgnwJYtgpzlIDmeJd4DTNqYn
kRCxLkhQUif8ds4WbsK6TX415hp01R1GczKEg9v2VEN4v4Tev1eLKXqh2Bs1gSfZqJrU74mligz5
mSnj/+uM2yY1mCQyWZUT6vZ8blECmWedhLwNH884Phj9ubEaVUCMyI1M7WMJfELRsFeypcbhwgtr
xjaNTJUmoflBzFSk5rMehxeyxGzacT2r+KSbf7+N6Zfp6AEZ3BgT9PX67mqWAfJ7P+BUDK8Rl2sk
ONGEkIZ/2OVr1Fsh9ZEUVGuwd6TP1s1yp+s37yhpgIp6OREbK5qO0m2pBx/41h4mvG/KGxA3hwVB
yUgWsWTgp9voaDyfOB7EvRM58HEcR6YGddDxMUkIfm0DbtA8V1WIIaTxOPq+nuvyQnyRvzelZ6bf
uQvfeffzoFJ5KXNW0p8/y+gXkgJj3VEsw+iz7Zab7/vzf6U08FpIp09JzeEjYtsBkDGN0+W48OJc
lvqdPCBZpBP51MKO0O8RMZn46N8dVrdVATUlsVL/vgF4/6SxUwE804lLDiklhttGjUVYtkBRZIAz
okNij/YO6WW86ZpWiPFvERPNymcevKoew/ZukhGUasYd5xsufaFwvzusR9UHv5omY7XVckxKjiZ2
n2lW9dpB6f7TVF9QdlpfbNp4mXpOP2f6QIVoTvkJR8kOrjm6MWr02lIc7BgJzdO2uxsd/xeTMNzv
p/UL8vxjFq0CARI1dnMdJEQzIxjK0cKrpDvVoZ8avVBK3zXWjQXvh/0aGchbxwoM2d+nylXLntCZ
VNpIlBAG+XNa69K00AfJlq3OSozWNrFBSU5RNMEbMdduRxhH8fpa0F0TqXd2EotVVGmLUmOYUx5w
XoW6mIbY0cPeGh8c5uvFcyJGyTofIohpao+NHPbpAgW4tHkxmW/VeKOOKq/otweCUOZVtEANMCg7
Mk003O7WxEXF8ZBJpZxhY+eIPbFXp45TMP8JvKwqQDvPTLC96XwziZhRFReIC1+IM5TyvcEBDy5r
75RTP+HHU2ne8ZCOtqZqnI+LiK7jZtWk+NVOAWgwpADlPFRFcTea0fvWBmpEvwALhGVd+Lecv+K7
Z5ioapNJvspC4+fsn6v6yieL1xQgw+hYm6+3AFirQSfOj+A2Cds6dXxuzjBmQ+hYAra6LAH6OkMX
SqivhQlF1R6JY9ER1DVkS6WPZZnlSqH4TgzQKhHpcBEscwh1DwXYZIEjYu4E6G1Dp70kNppDEGAL
wzfESI5tjUfe9zso/dcfv1slzii5EtOpOZVa0opaZQTXjdvSUcqkxJsVh6pdVU7xM1HAdrO7SbeQ
GwW1E5+Wl7IsPBaGxK6PPKheCerpT4hbDGBKmelybrVYz+yn9Loyk8FXA2btuBg1qzzvyyytv5Z0
a2TcUpC3nsey6XqrghZV8NUrMo0mLg1hUSuOSD1/wts1stYBvtCadRmycxlp2j5G4tEhGJd/+1XZ
dOasSH1x7esu8vN0hqdnut8lunS/meMQh+NU231OYyiq0fGY7lg0xBh+WEeVO7bD1vpe5mSVemw2
2qkIa/pGLD5ltfHq5lzeHAbc5ysXO02nEBtFeS0RNwz41B6+E00QAn5KfGkH7wj1UK/KjIJ5Tk/0
8TRGWPRYwJoLd++JkZGYabAIwIcRKagQoLYLxyyfUmBUDI5zkjBOOoYAVZ6TgheVTG2YXmj8GgD7
4ujDiI1w1hwkoXA12wHDfmor52EtrY+qKfP0gnNAiZtBIuxktE0ioHyLM4rHfy/vEEXtISIs7dsS
whq+fR0a0OqCr7Zt99vP6rf7zV6BhasIWj3XT9mwD6zOFjk8y9X7v0yyP2bbgHENyy8z9bc9cNVF
lQ4W3FTAMLngXlr239N9qwQ5iQUl7+C9G7A7vVFaFDFgvnWwVhTsaPpk6KUEgbXDuT9k/hVu/Us+
CGw8hT+0YMiLmpIgXGSF9MmhBU14XONCb080vDrkXojqM1KtHATm+ry5j5T8SeQoL0RbTN9i2m/G
XdxFvlum07rk4EpFMLGiVx1u9hvGuWhxgO9mgeMm+arWcZaiaHyfMiPpYgdj24c9f6+H9ZuNaGfo
1luRmRZI3Bqennz5vkK3R0qvlNT9VNynyFAvNmKBwczyTiCi/d8X2zmRPchIdSQ0tzDSVEGHN/GJ
1AleMCJXCYXOuMED9O1R5VXGasJSJ2LEjFZTkDm4xWNWAMIjaq8ddHTkgYfm9uuSuUNhbPkYFsJh
9hpaOF0WtC5b2NXdnjdToQemkRMYGzdbsH6LSAGYZj1P2RJ3/WxHKNJ0iQPTKNXjTH46kyf+A/5H
67furEOgqOgYnhNiSKVqdSU+50eBDLw/HdUIhJBkN5m56UWWf9DpflnAj/yKzN1k/E0ywoTx06Zq
J6u6z5dbj/3y8Q54eJn+rraudlTDU5XlSfbInaPL35M6yzfYyytKjWMoMS2CKs6YbZqd1F7OAwjp
2jXEiqqMV8mAnF1A3AT7/wcgeaii519ioSozP98+CUwMTk7xRY62m1aVQoQjNGKSta8IMaNlT0CS
sZvNZ3+uZZbB+pyqw5DDR9TFXacbMaQ0f5pvCfDhDxzFFJ9sgUowUzqLFO6ADIoM3hlXUOFT2eog
hNLYamkylOcY1nT0b5p3LOvF369ww7Z27J7g44rXD4mViBlmYSnIgwIOygzuhqxuYXAoHCCqpluz
+EHzhyBTZT0F20HwNpW9X9LSN7E24M4sto/bgnEORs6nLG5Ce1MXHgBpN7SW2etUqTGVx7LzIyrg
O94hCOsaUg6YPuWOCuboo2MWaVQFTXfyCF2+sVnhHrkt1VjdXUsUeIzoHHtcZcwDfxKpwe6TIFff
wnlgnVX7eh56U8FXfFM+otEt3zqqRH6biBvIzEjj6pU32FXm8ugPMtYAIzz8W0bEw5KTHZMNgC2X
4nNvr5RsLDQCQ673JYFUHaL7HoPGXZPJ7Y06rSf3hnKfj4j4SZEH/TmuZ3YywTUyxoeBmzcLRtfP
JPo9IS9gdcBjwAuyqAB6DnNwROOZguGyvc1j+Hx5mCOfXeV01Kc7DfPoXmBUIqBraEeTQzN4twkY
G/IdJ1jqQcXLYuXOQVpn0MH7OhLvrwNi1au69WzShZG+e4wrRV9lHaeQ4KjX3GaureDjgHyw09Zm
ra0sfrAVGT6fK6UnejErMEO8ciea92s74gJnu6692few9dhCs6tKZbiVf49KLTrtHqnK5RUknyID
VMOZxFjSOys/361XbyFqGLy2sPyAtr7XrOHgx4fcGMgouxcPllll23peGJ71B0GrLj2/R2iNlk7E
yNA6LbA/gDRj154Wa5dfT7jyEpqHj0Zrd9J3LuFDDusU95pH4wcFtfAv2MANchNL2PkT4pZwFJOi
YqIgtBdtxT7NiBsPCLyFx02AOpcMz5E9BU3fApiytq0Z9g89jDxSPQgKGipL0K8MfqFw3QnA1etS
Q0VLxf4XqDv8ZtZxtlPT8Gmjry6JqKnhOUsFLHyYfEeXOQ2UxCftLYnmUufUhydO7TUFfqcpFnkB
QIUonDWSMQz3ivsWJ9rpBhaBjiSdytJHTYtPYdXY0f0Ar1FrZsjWXipY06BYUw42AjBHpOpNkjCb
/KzHHtqSsPHzq6wzVKNcoCOLQ36ica55X0FqhMH5qKPXp/GavJ5zk6+bsaBf0ZX3aAAZ/kfvsK6t
bnDh85dzRDTTbvdBuxBrELCLHD/g10i1amW7ng02BwmuWRvp9uyE+RyU1UozmW1/WJQfqvGiR3cW
Nr9DKoHIWecoEmLpdMDU8E9BZHJldOtxO0diBL295ON1nhok4RXjWmstFpA3PZReHWukugOqc/yn
8CgcwnEQwIwjxBfIF7mA/v62qqfPenfr3TrSj/VRhplN7NH+IexdcdVXxQA4xLCpL+MjbdXDNNMO
eB18UMg86ksf7nOKxutdR90R9mIljkA7euOT8L3fboiEFqnynL0txPk3A42EP6sYYvDhHUlz1FaV
6b2G/hyi6D3uMvQV3K4AOCeeSQbXvHwS9eOebiTwgFC+1/HPE8wTughYIyu9SZUUNQZGGnAiILzd
10XX12d05CpytyppMydschXMux/0YAh/2Gtl/yHrM60E9iJEFb6732Qr3tpKtBXVM7EpuT8QcSsn
d2VJVc4+QEaLqIPzTkidvwRk1kQ+Qqdqcszxjdp9t6Ul71S1zw4mYuEeL9eiLWUzILc/uXmOGimE
DYF9tXzWPjghcK4liYxtK56euVFGtdYPws2PiI0iaQXSLdCHnjN1tYuo67WNAIze+YoUoI6R+oZH
lXTkW6RdxoZUYZwAF4IB0i9vIlhAfY0uWKJDuPZ1SQfRywVoYS5LMp35rVXM8XASOoDSjXTyCURz
+Q2TWYIWiJu+p0S/J6vOxKyJrhjhK74Z1UWTqoMehyW0XpQUralv3PSwhrTcoUU+yqw//ePf9Xss
qoEl7WT4qfGshRjhMnqfyv/dp3Oel+twvvTBGMlZO5bsjsIgMqvjqB2hJwV4L/Q/3acoDHncsaep
+eb8r96s73dDSxAa+khIrXDD0QGEO1ECkyx5uekGmrgBTHHGywe/W1vHWRpwfnWABHTGw1TmHbYY
UBZOsVqDBB4uuPYgi+wuNLmiOSFQxwEEfC5a7ZSkP44XfIVuSEtSzewU5HlSQq0qdiBzvar178f4
fqFP2Pa7bbRWazUw2HLeV+zY1ORY0QFQP9ZzhNVyzmrXf+FobOezkZPJZDEMK1rYUXkpiYAlmDoF
hDC4xeI6nP5JWLhzMpnKkjR0shIq11R1O8YVbU41DdSVixysjhueoF7GIuJd6kkSgDCDfHhItwdl
HoIpLr+yFyXO9Pswy2AQz6GN779apCFTWOyqbj2dPI1YgQkwtc/b4QyrIwMuso6tt5Evli/dhlci
5aBhTTvcDUrWPK87UWZDe9LsmScOkZjkvBJG/k6cLae4loOSDvF0uf/oKz4tOTDCWNQ5uBz1DmB3
GJXxAjmT9cOhh2govkY4ASM7PGjRlqa6EsbH6dNs6PxrfaIqqoNdAEXNnKehjHdzE//zNrYXE532
MI/smci+i2Zoqd4J4EvagtOjZfm5La5MlYzdNJ2rAStYwIkMj5oaqXBMAcSJBMHHebVxbePMh1Hh
uxk2szEHZM9n1aa45z1TPnIUL595m1BdgWP4B5UiaPuYLsADRF7uLjCIKq9VCN4n5x84c1Ug/kKd
S93HERXX4KPqJfHXlU+Ts53Wb99X4KTf+vygtXFRA0Ro5HOSGB6ZwD3gYolXkobMs/JQnQlWboro
Act/u52KKz6CFpVc1/mavvr7TCc7cO56OHMBA8pwo7CQkldZ5vJcVukTsPLsKMBdE5UL/gvaRQlO
vAb5B7auyIWswL9uSDx6EDC90PqjKQX/JibVtPH+rHK6Le/AiUWimiK0XAndwitMHDacABZe55LF
AJn+ybyaPvOqQqoVx/gvw7x0FakfI5gPO4d3diJbXoZUOw2+hwNaazU02amh572WqrKE/BZlXBoe
1u5ix9xgTfSaz5S2rjE2xEe2UrfpgasmxSL2MUGSuMSSIuSHtBEUm2fQwgODkOqVa0lok3C2FHJP
PHKDbM39S7lr8wcJbMm2VznYHqzFf9cVglqs4hM7CzcgKQ2zlFYswrR8QMcxnRNzQ5U+JOVgmQzQ
cyyfY0sZsEbF5ZKkAXyX+LauNsdAtax8UFemA4vOyMkyhqZdWqJdQ/knXJMxCZ4vhGDEVsHXP1uS
8yVULIjHzbRW6MACJjgA8V0+hnOiuFV8vBmyy9ztgwuwFKxcYrnYjHdUoxrSjjQ13Tpslbvdk4I3
1TEF/YMH9FgmkClwcEqre+na9zhFMjhikxO+fkl6fDRu5+wTe1ItV1xNoHTiMsDgrexpC75eoqrF
ZW21r9djDyVhqeWHhyk1xg2CZVrnN79jNlhbo8E9o7oX2BgzTs7oryp/DFxpgbERtTGUAU908ADF
IjgNlWhlbkvZHto9EF4HRJ7AEi/km872UtK0DlYWW/KwSa6+0eqDQoMWXmsDUqrFXPKaZf+kUwPT
3vz4hp1tvaZ7sbYZusMSpAqR3DHKtPhA/eHYyb0luyI7mXNI6XBEx2hMuWLoGbcP+TYnyWM9EeP1
ATPSpWELM3hqQ6CD6TSI21+XHxyAo4m/uyTUjAQgSsxThe/BzJ5+xqwRLIgY85HN5qrUYz/QX4xv
nYzyuSynvsfINrrq3rg90iYa4+gbcjHf4WEiNuqyM8TDSv/X6BMsR0WBmBg1b1LePzDZy+hPpfFG
+zXONbJebktN02ZX1cUA9FOv+ij4t0VRbb/AvIiNZUdhDMeegg9tCtkmJp7Pwhi8XvP13jt1uGcZ
UuYHeNoPeKzPyZmlJ+WQ1onZBchPiEJHVaZN7uQiu9j3KF31WrvO2eq1qSSML2KOl2T0ecnJQSck
iVevAdYjKzizm9hascdU9GGXo3USD7IJ6slpVzJS+vvTZLV0hJEJk98q6qeaXO5rx4sgHwH+x9T4
G6Ko+vRVfdv8wB92pPv8oH15yHUhYXqmZMWdVH5+RCvd3XxwKuwXydMqaTePAgSs1IHbiOYeBGpi
2HkRAap6RDvP39ZQumw7W8RZDZf6RjF1TH3Rg4l1LE2VLLe9fqRrQIRVf3jQHghbdplfbjWvIWgy
S7vayBbCkyRYqQ2+5nKLRMeppN+QG8E2swMEujVSG4lr0olbxYCHDR6+nGmcTq3fiBsw/DlZIdSD
/u5Hze5kfyVomjTfzWaQDOlvw76IaBYc4Sft21i5gIxXwLg+yOsfsHxD86HhR1F4qWvvGQmXEAVd
YvfOGMsqV0gNbDLoQYjQDBrSe53YR6koQZ92bdxG9SWFs99hPUsGy/ANrDcVrSBMYq1jSRIbXGDH
SzekFdhFwjtTRptfDrkwJQArl+MsKWVaSu9e9YMuaOOjNrFkRdNAkhIxXwI2pxOTY6T7D3MVd9HB
UbzOkUA/uBfZfLgx9IxHcyYS3mcbxPlseG1xwmUTJOGiKosmwEzHf9mb8Auyejd7ipjz5naN3CSB
4M6891ImJ9LtgWk7LhYZpDPcWnZNh+kr5+1uhyrUvdMlwYEDzMC0NVODOjjksKAY8nJEy2q9YI+q
fFo/GhfWinu7hvFMfTuC71r398z5MJxj2RBxQ7EUoG5LXHTuN5cf0yZmxuIMTcxjaCf7spuJJ8uj
+E14XGe8GI1eAgNEzgIoERA1XMPBjwBCkuQxAaVOj2intiKdui0q6w05Fp49koEFt+L/6/U/aszV
5fIA3qGUXjQL3IYYo7t9MMlt1Y/rKF36iXsNjl6CbFW4AR3u2MA7liVZuA5j1H6mPRyjwYzQEony
XykWyEmbckOd3uI/Qgm5mcIjUdzHwtxuFqvuA8W6RmF0Lfy1Hv7edpuAVkDpO56X2/wRSnWKg3uy
KWnCZvwIgqS+oKXYpur1kCFkAMTAXQFPbQgt3MGP9E9941TmkKbj66wn0my52Rhw/oggI0019sZL
2WKWSLjVNRWj6shO/62py5SIZFhaWvSVXqOKMsQy5QW1HcNE0FTGwm8Bs5VMiNAsVv2YQTmeGVak
VPDIl+K4ZR6e3MXRqbR8LgA2q9783zEWcnHkaTH47i1Icvepfz9l8/08Q6sPWE+adVURvBIzFE0N
OPNuN7nKfyF2l6Ab8+QiEUaHhXCoPRDd/A4cNl0YvR+oBbMyoGJEC2opuoiz83l8ne0Umu4FTN41
Dk/WHWtgS/j90w25grtJ0jS963bxylgtwqeeUllBxKAq40Y1MztGSFKiwFaHQMOEPRBbtLyNJB2I
0+Q52vri/WqlmD/PdutOAHUqdgnw1e2/Czhq1B+0DPsKUkFkm+s50kkFZEyihs9PgpREWtSTSxA2
2CVCc5jIaY2cn3QOO2rjEFdV337DO05dIqvtai2kI/16qgbtY6JwahDMuhZB1scT+7qkoJlWPU/D
D0D4GK/k7F7Xnh+/8/9tOZ596OgMXmfIO5+33E4seQkZchKyMTTC5pkbTMhDLfYTq2pgF4dX6idX
CBZR08qdTAG3ufbr0fReJE2NB8oym5fwxMa58FXSPGma54jN3lrMzKq7YErelrhzFEZVU/qC3avX
EyNJ1Ad9F8PIkzhT7kBiIZ7yd/r7/6qS+LxDPI/0EQRf2wJaqMkBGAxS3blW1O1GStNDcGAZh7yc
MCSbBHb4uI1eW32w88oZecW3XGS9e2vLZqivQgqfFCBu1IeWMjWToKOeDVQdWBTGwA9XpBCq7vsU
NZzCTyaPAImSpTg+2NVIRF0PT2dlKT8US+VkJbcb1UTbEzkT5+FsT+6p1sJWMOepB+Dwd/9qdMkL
sEQj1pKHf2+ELwa1IB2LwRbb2yhbM/bTFOiSrxCHYQQkUgYEJAJzZPpMop1Rj3tkDJoYFNAxn7W3
zwJJ34nIRNvhF21cHG/BFcdhs6pTNArrAmt2nyzlhyGwbP5xDorUVwWlASNMIWUAD/RtZLzE9khO
zJDFxG4i3kgnqWKnPyR9K4+dv57ILebyJ+fjRYX0hPf29y2BiAlqygR+F+axbe4ozEu6pGHwGIor
4KFOdezUIzXokw1XcExiy3apsisClrjXK0Ro8/oKnClVe5mCj2LTAH+mwl51jH9qVH/hvfVCtruo
4wE5RrMxEm7b+riPCu1wHKiSj+gyzqwIUOoLbJCohxiVI/AAp95X/3z3///RDlAUweqedOS91UnP
Jhsn+jVuA/xGCfSMwK87M1dIcrbEACx1E85gvQlJsMgb4CX2MZd+Y12Kn09S5xR0zPQc+u1Xk4Ig
nbVOoh3HuPbR8Gez+qWz/XG1/VO5VWVDPogHR6sQHee/9tIsSRdc13ADhkAqmV5M8C9iFs/nwNS8
9wyh+AOme4w6LwLVoF5wLypx9vh6EtEA6fBQ9+37hNE1mmCMCnb2Al1oyxY61FV5q6tY0t3/iGUJ
tnJZi9IassPSZPQ+mw3Qa658jBtybSNZGpevcg+xLQ76fK7ofU8sG3DgplYu0eZwSR0iojKU7aJX
vuIbrsupacDu10Spms73W+igztXvUvJ9VKypKJL7rJIONqpgMQEvcWb3+7x5Gk2V43YzPpWvpK1r
gula06pcEmRYdk3cG8sthI3uvAgpraHy+0juaO2NAcodWsFrHDOWYEFU8OPihUVbhQE+DMrQ1Sm6
8tQTK8xFh/xUWFwrmS/5mAwCRDBu+3wZKxL0r/BGFnM0C1WioqRbDxeQwsDkxuamDiRdYMD/73U3
QWcdziEtV/ueY0CRObdFmM3+iaUTjYxGka+BM/bJ86n6tYew231V5iYqZP/hvNfH8i8P8MP4Izm3
HfOXUNI09Neq/HpxD45nKTA1fnvUGI6QulTRpDTQzlw5fBvQ+bzmRKv8MT91yhDUqGklmnoI8wG4
O3EDahsMJqBT6Tcp8b2LLxUiChFXazVQ0HJleLGCjFQ2oL6WTJ6EqhgIQ0/0S6LkmB3AnMx4UquI
nEKZHoqpf2OpXJT+sW9R2/gJNtDQGGrD9zgjaX3/vPeXDoxhPjJ9pGGJFuIfL7H2bdlrn13neDE3
BItN12wFDQMhESMlpkLmfp2Gk/FUxqxjzfTVXuobMvfrUZRkZD3h44PJ5gyXFvnue6jqti9S+RQK
o9QzVTCaKyO306Fyeyy5ay/0mBqWPSlkPBaqIOrdPiSheNvn1W1Ij4cxgAlUN+m5pLmbYHc5WLkZ
b9UspFgGcPHg4a/u9cr2xQ52WSoBYq1v24bL+iyJHjc5Rum1PX5AzOt+NuiazOI90N0IqTgwoUMN
uwVKUfOeGi4UTaADHtd92Jnh9qkkAYmUpEDk8aGwp568wNZ4ut24tdRuGq/48Lq9u9Ky3wmcMC4H
G6JgXAz2gYVvnJD0qQiqMlhgHXW8JT34XcT9PzZwAhS0kLKDmbYZjVckBQ+kg6KI6cAXYpHcC6oh
SXDT9kO0REsycq9NC0NBdh5/Kk9wLMqoIHrxGbkMID/DBKrR4GKflxnrhab8CSNbqq9cXQGjYHlV
3ib0Qak+iVZ7VPap8nthq95HOtZl/aabE5/Las19hV6o35TvPd4w+pZEHVq3YpTDfJfxjMUUn4CS
+WYYb3Qb2U1zbcDqQh8S6wH74C3je9VXUEHA5GPTXLlbmNU8ezkr9dVRDsLhiUC9fG3PbWomDZl+
ANDFnQAsDs/wa8m62gWQPks6M0OCTlxe4xO8/weZ0NlkLgvnGDxzQyfenqVsgNxMpIrRWG2HVoA5
TVxmG+RWgE+aN9Sp6FzlowJrRSRL2owEtiDJMWO/T/Ny4FMwoDfiixCoMFc8HzDuGnw8rjuIKynD
GOQaq+yXjOaZ5+g92BhYPg5ZsWXHZdF2DYfe+u2k4XP1KrGT5ICOGREvsuYQhRXySti48Vp5mm3d
WpfQHk3FqBc743ZWlSjLH7x2DK28Hhy7hhENjepUdvcaF5xH42TjdUHaj/GXvt8Ec+9WTBiZIZrE
3TyzGX82zbSCs9m3glbeqFmxpTpVZgUXRyTPAo5jr6AQNGA9rP2O946WU6VitZVJeQK4wPdZq6R3
HAcbJ7YsI9lRuYCOs/dCZJQWRsl2ZPoFg3My5mrf5jdktA205YSaQvs58JtsHY801EpXcGncxFXL
TiafNfUOCWPgvhBjqwoblXlg/vTPlY628jIIASG9gLGYE6g2WECr6qh4K0iLv8MnL2yrbm74Inyx
6WtdAHKRBm4+8d8ee2M4G1ntpgMxidasRo+DuEnMI5UlgSu4Zuax/x7m4eyETA9HKhKm2GwOiHPZ
FhXMj1DOKFSLCk4x3GHJUn+VcmmFNnLQdBJPaKk33PbR+GJ40HYw7HHzPvFNoXwTMpR2S+LI+4tA
djHs05NexmPa5apRBD/PCPZdiaejszppY3RJe7N9SFL3qkxlrFICOj/GNHUi7Hdy1k7G6QugaRT9
tKMcA416O5HOe4iaFIcIj50DGsMfoCMXoMMjaYcWomdWJIoavxWajkfH/+7EpGsWhQQikahDL+Qe
eleLNNXN/cF7zLzXQHIG92fzsxgZ1PrXEemvoIb+zKBudFsQoVEad5NeeNZSe79GzMvdlB/1eRRB
Rq6BTfQU9HSWMqNSHHyWVz3g8VexeZoLz+16TVPbqK2372Ea2BRZPYqa91A4gRa2ZU1du2qgRYnu
jmXjNsRljlAybI7Lx+DHt5UJc+bqbppzVlO5cstq0B4GE5kJet9nj9KR/+Ehqd4SoBj4rrMUZEuj
lqdqan5eh6/SpVhxBQChBYPVsz7rCHVLM9o6rRP32R0qnlGofz/iyUy48x5qrKArbpjxJzymumMe
wd44x3IzgMepttjJDqwdNpCOEzOHt+dUBNre9Tc5gVlJJJBWGBkX3RVzHxzS5Aga1FrrqIYZrn4H
UlrkLNHLr7ny7kjB6iNkezGBWOu2GFziAPH5bbVQztU09yq4obpelmfwZHlDtF2NlM39Gf7gsnYI
NOFlYvPn4jrc/q350Lc6OmJ0uAXvgJNGv7cPrddEov0O0fiPh/2e0X7jROGUucorjKsSHK7Q7qtn
AhX20TayVaPjSd66BUO110m1jOFKlG+0Jif+OQXctbJdQhjQ4Ix4mJtrppzTIGOoemGMJDkPmWWj
iLKEl2QsGLsNSoV+J7FZh1VkpiwhFl15upPc21ggMGxwWg0t0R8HEpoL3yfsC1AXCFwTo+xe/fXX
9gEjIiMWqhzKHqHqDPJ/gaZe8OHT6qA+yqTOu6wGiww7RrJxTKbooUk+2Lk3OALZSexXiUDcsUyL
fX1lHF2n5Mrb2f2KjVSxDpPucjtwWLVMVOb0DAz7u+pLwPRfLRtTuPAwsgNSxmVho+o685vRWhpe
CdJ3oLPYjmdQD1A1hfbUTYArhKVg8GfeEWY+MN2WoFKjPUF302gKWzmMUcVC43r3o6oXkEGKrIMn
SZ+UJwJ6y9WTvORsEoDIbX8hAf/y3ktwsNQw+Yn7Lzp2ES5ojii850oaAA48ssbXIOzCpmza14it
hkA4mteaSz1DbMMPL0d4GG0P6DjX6QcxOq7AQB9uHG6qZ86sU5YzqlqlwvEuzo1UILn7hMXG0oEd
ysIq2kX1IBdFWWuWGk04tR6S/2KkWIcgO/fVsgWSroAKa2X7cO8dJo03eb1RSAeORX+SdIO1nHf1
vDmmrig4NZerJn52Q/PSbZdl+lcUGSoJueN6uUA9NgqYNPBnZTHbyncMieEK0QhjahVq0ah59jQm
PWewheO9gFMD1sFvA6yL/VaAIDVdzDc71F8mGAk5YTYirSnhzpCAdEiTj862bojX3T/4Dyks4B0n
MFRfEzdWEllFR8yJm2lD5+E/yN28A5Gt0yXW2xsGXevtcqkKfEOoSMNyZsx1E47Xsmzbvj8NsfHr
ZzMkB89XsvcB3hQFIlWkzJvBSWLwSFFWQp7xy0lRARqVkjr5zYieP4e2iCm4MQeFOr3HNds+hMTC
1FMQ6UcBr+lNpJLAv2sQadXxMQ3WeU4bcKcezTRjmAhFvzUosfpzgS64vJstEse+qQx134prEpWf
J4jV1/H8yxnEvMBaMcQDXqi+fycVoP68fFwlLs28Qal08jVaU3qXmLjIUMtb697FgMShkdHaEbYX
ly6D1TiMKRef1rR02YqCHpd/olCJYsN7fkCAkHTSYQAORdl3tzqlR4vLaSe+KfyeFbGHDT5OG69K
ZzJCEYa/V2cYjemIQfwylKoGs2ScaPeuwSLAx39Bb07yD9xsQzOGt+qQ/0VbFPU1kAcdPV0ZXrSi
W4V3cqnAS4b71854pq80z+/SRoPugI7VCAkMdVfhTHW/NqeyG8gPZ/5Cc4l86Ql767a9N4ouFeHG
Gs0L0RdrHn7h1OxGnzPEhjn9P3LuKmO+SjJI1ESpV2TbO6/gUGkK4jhBfDQ0/8WI7G3BZCyPkiTz
5TttiKNv2K2GQdEM24RhdMPE6mVRyna9o5Oq1mQW4FWj8ExL0TFVzPostac/eOAYdj/huSXrgC3m
FBdWQmD6lGT3W7uw+HrVowPDvGcySRRlGkytOreMulfkH5S3Hn7hr5qmZW0kJv78uGKBDwwGY8I4
ZO9dQO3ShSs6C7yOP61uYytQkk/CGxLNLrOFsWvuOJ2URxjsY5jCo0mu3F8mA1PyvTOolBWWvsaA
lmXJ2oqtf9SwJEWbWnHvuHLtG+K1FkAF0dOH1mUErOCkp1sdusNk/fJedGIkLwV9a+xJ0L8rpNGi
nTcVdC1cGO9PxTwCzdRkP7f87PKdBhCugo+yg9UYQ5w1xrtdpJ1kh2OTkK4ZEuOGMxDmTh0QkW7D
SajBtyUSfeOmh077lWL156xILTTAYzZMzDLFw/SQ65UO5o4An3qxOgrUjRg6xn7OnkeHJj8fjJb+
ZesGx4cUDIoQ6W7FBCwDtcdj/mZBllO3FoK8OBF4tHPIROQUwwHtHjwN9fm2PweaKeMfTkYw82hZ
ifkGHQQCeHK6VEIv80hDwduGDyJFBRM8KV6ROdPxuUlF/+IuH7WfRsQYxh59iD/LqJl2rGYtQo6f
F3GM18L1m4muy3MFV7MebzEa62vOd12RmWQmuiUbNanmDYDiy93b1qiZe5+HJL3BdtPvT4nN5OEU
2v+OVLq52oQI95U4e+g0ioeDBPqd8byH746DAbv58gEZQCdWOYVWZGzdp2NRTWc1Ocxh5M5LHORp
5Wi4vT3DDTOAfY1sY/uqVWlm9phYrRl/xXDnxJllxyN0gEnj8cUM2ormudakreVKLlU0mYcCqKxF
gy2Tn3pn90TTP/9q7Z9xc1KOMokZkUDfoqctEu1YL7FdvXRPV2l97Rd8BPyJFeDaMGCelh9UV2jn
0zuWAz77gDKwvDFkLWyP6pZtblHGS4xJWq52f5QEe4+IAgldEKLI+X8YXpGJhz53mFZu0/cpyIn2
VmwNk/NIKvaKXinOK6yZsNEtP4vdZD101KxRrOz29Qij19TgfZBEVOEPcAeZcPXthRJFZD9wpXAj
9HRfrQDyg0arfPMvZM/Nv4xJzq+gvfXSugt8NeqoTqIM8VhNMLE8qAZ7CVniLs2+8Hu+Uw88MHqw
ioxbDLWHwb2sqSw4OT3ZK1gtmMLUsfBGqYs3ukitJ4ENwZC96Mxc8byXnUjJC8mQQxHzCQm++kC+
5KEhAkYQE+qqSXgETFSqT+bxTyq7ZFK4AZT9JOtVORtMahCkBnG1Hb85pPOYOk/BbWEm/LsLP92f
c6eEe2Cmte33LoRYYqPUIpZVapZ5X+NRCCjc5j0crPtzBpX1iaKLSH9QMckjk3jwOsfyHLavrVnH
7RoizmvHLEnUDJ/j02qSje/y7hp6bqX1z/xt/+WyekutZVa4BsqK4WcNmhdJOrwraTVP+5ay9QEf
CdJwvkzWWwHhCslVAdXlckobfCLMXUm0+NNFd9D3DEOo55ms+ikNUY+47iXTJVxxLamQgYnyAqQJ
/Pg8wHVQDEeeL3pfCO0Lym69D8dZcut2rTwbEmCYzfpe66ZNfmSPYdmFKwgZS5AZ75XwNQMwXuid
TSIiZ4P5Lk0LuNB9S07UDIbDhTSYkRG0Hx2oaoSfgPecpyJJXe9w5LOSx367nABUiCv8XDFKDx76
R0WLw8LoK8SJvc5Yv9PILRPuv0YvO/wdHMH2Meil/gvDATpvb+lHvgLPoQbTR2iLoJMgiJGXOMKV
p6iGRQXhG6WP/ja2mCHvZObQIqx9to1GF6P/GB42+cVynmg1LRPKkjCdV803Jikz0l3swTg+UJ5V
8Kf4FGm6+fwbVsFJu+HCDkBGdVJeUNWLA/R/B+bv+KqhoOcaQLElwy10cKjLMkQ5K28RMeVsoAN+
iNb6KLpqyOHiK4iWW8tlW8ARzGyxpaaEf7DjAqt6Zm4KED1H5RmnUFbY1b6L+aJ7sxYzq2XZp7Iv
DLVEo2PxyfSAubTnkhId5XWC7eWlCbGlVoRKp1bzY59pol1s7d3YPzTDudkH+XYR2jcPR1CiYI1/
95N4x6kurgB5V7L9ZrTXoDS4ED9OnH6fgOhky8O9+eUrDiybDvOxGHOTCKRmP/xE8ZcR5EWYN1y4
8FC6TtP/6diutcWKcrT12YI51P3ztubNIHpP5f9bcZAGRaCZveVi3rc2BBhkQCkE48Wg6TwJ3aAv
LEnj+kafx1XA6v40Vy02bwb34pgjb/Fe/3OoTbEBpMVibLvOLHtS507w7x01hzydYkIoBHyx8dyd
3lZftpiGb4XReJH9nEMeQ6ppcNeuOUUPepds4my8Q4dmLo0hp8W40zEfVTPdRsPwAT2DgdejAed2
e8nv9y79duPZ4wogFEEwrBG4L9evgX+AiyDjmqygqrzdZjcvFHb4aX4UoFb32fpKjyUtIdnhbZin
sWSyPL41iM3B8xNmRoUGHjiniLZIPg4bm2T4woMEdBXfJG9RI5Jk0NFhA6VK73B4axSVUNnsQhXK
KXdfSwv9RTYpMfVsC8IF6IX7sR6OqGXxtWDaVzJrxWvFtm+tmTNrMpr05UDb4lTRkI7T8IQ79jGr
SrDbjqf5jjm8QoN8hdDojg/V7SFQJ3ZSCPc5sfts/Qvnj6ejkl9qbQSCroeQu5+g38KC93Ccm3hA
r/91O4crbsCVhwjyFxhaEeeyCQQun39UWsT2jqiPZAJCzO0nQHRo5FIiY2Nk/27qZHwh2yw5UWcU
UibViGta2Bu41QSCL+BwVsg2n9/OzDxB+Vkv0MqX6Smr0ARSKehs9Ogtx7ydwOFiXQkOiPmMmxU/
MSYQnC9rTuQCnKVgH7QgbdaEldrLfA35CqM2si+fvTeodAEunxx/jw5s33FTcIOX4/sfwHLQ/MRM
DXYlxmphfAARwsg8yrziWQBug3in0IadkVjqog+4HbIdFNZoeZLAGDrIeau3ElyVbE7LKmpkxpWE
j/RGLUIQY+UB57Bff4XmzoVBx+hENEjJ6UEAaApxnzTxJ0VAYcZQAce08XCI/KVWeUqBHMrrvCm5
/Upsbou09WddmFTm2QtPt4IJO7HgkzGs0MtR4xLkBAuXvXErGTVUfqv8gc4/tNfhuWKirf2griKB
XHpuJ83FVpN+D/HdBgFcl5y3a+HbLw4M1X889pZVGSb0DaVkPB8XBXRn4nlNorCHCWD8EzDqaDwh
AliJ4+RG4cRbzSoaP+wnHF9QogYnEGwzrCr4410R8o1eZ43WlDEvcmh5u8azHK2Jrezxhp3gIS0k
1SWu1CcuMdnwCLkcXGLgAV22DzzD/QxW/WcwIdAwJdDQ222+NBO4UA3m2HPTeK2VeAdPLdSsHkAc
vHPsQsx5To+W3aRfMlIeTft1EFKfAe05wZKbqQUImjnQGvIk1+b1S370Z/aqOzEqkhuNLnGe0AYv
KQ/cPKmUyIGowBgwSOwpO8ZRi8MaFmsmGFgg6rZgnLF9xO/9ej0tjSalq+5ZpCFvwtQeXP/rKEah
p0AGChrMx0XfmhPNnRnm9zYL6FCxwB7jC4pA7pOo+y9kpY1yZkzHTbBIwpmGpjdHSejwikyE4SxH
z1hrtZ4O7IBi1LovltL3pAcY0U7F0x4x8Gyoco+AvFsyFowBeWFCeybmZBNRzJeOWsyqHjOKC/IN
YDsNIHdbXMnojwpKCsW6JHUDNpyHYws+88JJjXbomQR9phLlMQc5vA4TzdPkxRkcwz8aTLGFNCGE
p1OnDJI6UYDbrcrlx1xVz/4b2vFFNln3fn9TnxuyitoExzJzxw17WneVlrCcMlpfYyzRvwDE45jA
IJ9gIhxE5RLlybiA7df8CBVw8kS5uOQUylfM8rZ89iuwS7CyFRrZetLgCro4qFJAyFxhon+MiGje
vBmE7kr3+jiAZ66hRiT6r8mkxhoJ8iUVTXqIcMbZed/o6OyxUUtuGnMjPNuiRC2ER9Rk9ciuPrPN
Kva8qnLMQRf5r+WO6iWUp3+D03VBu8ZqK4vC6GQXqSe2d5QbVAFYo2iHj7liOaLrIbXI0W2khGNb
WqAGkOEBw8+RUIMFlgkzEwDPKe6cUa6OybdzFMQ9K/dOgZf5kG+V5pGxAhU35irntQaNehkDRoxB
oH+sZ98kOMa8ca7J4p8n59WKV2m+tqL8rBLCtZADGNIUlScogIcsnKQDRap89MXQNQbM0c47szmL
temxgS2adI0tvBRAqHDgRzO6oO1Og6BTHo5vAwsKXsyS4mATlZEGqEh/+76I9ClCs76AwEgVB+0r
t2JCeCSbPxH/6vEObqyKvdvpYLSE5DC/6b6R0OXBmiKVf+TR+yxuC2frV0LUDg8Do/OZli/E+WWL
tQU7wntD2e1IUnWUg52mqdsU5mLBFSknZvGlvUL0hcmxYGopcvpXbWbU+FOBkw8UZye3OxoT92vG
swkPeETZnrLioU1zka2RenrvkwJe83AUSSIjNGuRp8sIo2Adth/QXU2BRF2lhg8higo7EgBEPGL4
xQtZcbiq3HzAyTv43MO4mdOq7xKaiW/VbnAQEz0ZKp/PbUBVomel5h56rll++ylfQcFpvJpMl35y
cP+zkpUDKwt52Fo0G8EYxV9xbjCLNn+gs6gYAkXV8mQE47mBuemlroGnnRziW2r+1NijT1QQStk8
z7JiFdhHzU5iR+Ic8vcyQoI+ReSfhQHHGzPeK6eSGiU4gF4B3hKgEdqnYlJfZnaYurnp/RVHlh+E
WjG+6WW2sf9KaA7Iq7xFMViclXcKbw1lIi1wMzi8J2hr+BCTIRv1AGbmoK14ywGMBuXiTAoeqWrU
4mBV5jFydyV8hDMJZLb7lNX0aMv3PYIp92Ya3boiHPLdQ9lrB3WdYt2HJN/wvFU1F2YCstvKUilG
iRi1ykrCVoNWVhIyM6lrqo6QWYGSjPU83m6mg61Xu9VIiO4KOhfvcVQZ3BEuV+Q6p9+RqoL5HTua
GLDeTsCaW4BqOzZnIiGh5OeOandkiQFVoOz7VxFDCqwuZ0Oa+0z9eKouDBMOgokGgM2TsX9AO798
IJB8hnlxSC+U11GCQibCP7Zt7ZzjskQRL6dsEKj5fX6EyA+lE9bKptUSZRJ0COHg5QAyXvxD5bI7
v+6bW2iqhmcTcyflzc7eOPvnV+ev+IQdyDaqbteErOtYpIx5LJ3Tqv/iniNUOKaqlSFc2xhBAmKw
q/lwX30SOmA9ZLwgYL2ZT8hbpsZKaZKDkRvE/BYVehz7/Ls4np4vxoqebB3MUHaqs1MckbATfxUy
2DxLoJttAP6aG1XFqU0a4SiXntig/TNPi7/N6lL0F3Hza0LCiHL6RNOP5z19gsdpvQvCXa0hx1A1
ifUs+pSf+bqXiQspQPFLLbcZ69CLw67NitwdyFejzStbE+epCOei/E3ma0TmBrVVOZ7+qodK8y0q
p21fcgjIEbVXgNQ+EzfuUza0E2UVi0/NTmsTTar8+AUG/8IFy2fscVkE57Wbr6YbqjKqnq33o97s
pZjvovmVj9zMqLqU7o7rgIn+P44M0V4/LYW7G3gfcI58QUTOlncnt4WwvkckEtFfEoaNvfor5SD5
K7yLOrVHfZYRGn/g8hiwyWaULOWNe7PkVxJ1Hbik6p67sToXDH9jZCf2B+cFoaewL3hGP8Xb3Paw
yug2T8lwQ9qXJfWXU7TWiAXhucqICBqYiArZUjj07Fv3vMvHD6yJ+69dfRKbQbuA8A0qaz1PJZsd
ltYVXW0ogCSCQNoi44awo5WOmar5XVdy0yZRx+QQEZ6X/qtxS/fqboclIx2jqdoFp5kPJ/Xr5Zxh
gRDVut5TSXyjBngN6yRhiLHZp67N3HMv+84OJYXGEdMxk8EpybaAnpuiGOVNX0sIcznq3fx1kMu0
Oi+yCOBqs0/UrMhWYB0PYhTjSSwN8Vte/jWjzugEdHZwhoKrprwA1mzdNk9O/SR7N/Yen2j5Vvdr
dhhj4IqN0hMtuj/hfdAGUDCG8B98j7KVEuYejEQfzbgwZ/+zzgX5SthkJnGVpsNGpvlrdaBFy3b3
GNHLhEfyYAOERSAwVaB8ZbG0Sd+Z0Tw63u08JBYgYDOVlB/rlDElS2WBtzdysnL7mlHhltcYlHAi
mlqJ48tX43UKoxW2KpT+HupEVYAduvuD0d0IZ8MYWKVhxQ11UuC9GqGfhWPb/CECjok4QAjW6mcC
gt0vpGm6z48FLHC7gpdkBkjSgwNMQjS72kfKRXceOZtJVlLa83ThLdgJYHAwpSc6tmVWNbdfRNMb
0dPMvF03vcBegF+1tSpRK3ucD1k7qLRx7OICYbg1/eh8brPGmPXCzfoXx4FlBt/99fuwmxjFAjDw
bQoPEd8fF1XrKFgfF0ZXuveiYKFEWLz00MKSpUzYNp8epiDWIOr1OuxSKJO1AE+TpdJkvP8o4fwO
zCJYRB3YWxkf2ev8n4qUiu77qMtgt6QZOeWmAjCSs9fDFrwKKsNa99WjV5SpvOTx1TZpRCFbzC50
5IcyeOCUjOhShIS5PxR7lsQ5TC2EQ7KeE8DlwUKciByxoCARmmW8xMPYpaLkwZ96EQVVWE21SpQO
+D+5oNPurTBjCdSXGZILxY7oVf5UnN/XcQBbnW4gjs7oH8MzXyamLUVqZhWBI026Z/G21CTOYdB4
RvfUdH8OgNhzS1XSP22ct+sFycGSBFHUBqzTL5kDI/itiMLSLiANMlpHNyHBaBgdxapqmxwjewUS
m+ftjc3foyGmPP0Ztr+q/+cAGSs6QSxduarzmOZxYnU4lWWs0nMKnGa0lPcbPoc588dYcRqtCT0i
AbkSYvL06pD8MoHW0rm/I+ujrc7s3YIxsGbc5vQTZf1ccHHHmGu6sDk7ZZo5wuffqEjjqN3H9QXK
v0pxEBjR+78saC7ARzWQi1deYerbbYCjT52Z/t6lCKwS/tJEnCmNNH1+9AE+ebwCMe9UKcwWC3ig
UOCOdgO3PP9Axk8S00ahDKirmCUCx0AKoP4VEzK3pw231RizhLDYqK6HQ6E0hk58yniUjzICYEy+
4uP4i28Vzz75aqI/suwgLj+ikJGrhMvWQ0SdxfHjPpjtmWT3mn7WrdTdDoRogXbMBxF5sepfkctM
N0ArZDY6tF6XNcLGV180gG/zrRN9vV91PxCmdx6elBfIe2H8NBq4v6PU8HwvX2O3Ow3EsbTw9Gyw
xuVgJFgTTlLepc1XByCgiVFbFqK5IgzxxpIQ6NEFgBKxdYqBfQJz6AiL2fjhLLBL7JxDHyiqqGhL
27SCtM2DR8x3aUL9EXwgNx7vDFaqdWhKBXrU+Q5PPKHgZqClNAjkggiRlEhzfuPYo5K+WnA9T49m
9etFh+vgkDLbEHhCVY5Cz+i1suEkqWjR+MFvCnS93XbI/YujYdjjM0BQLH6Tqbm1aqtZaQ8gprhM
R9FDUhhZ0Q05lf91Mr8e5Ge0K89NURtDMfDbakttqQm0EqzrxEH3IubYiMt6W0I/Sn7zcGQ1N53c
tUdCGonzUrbr9++CIiiQth4dBv10LJo8qZCYljyFqU3XY62F7N5UIODAdbscVGEjZxdprmeQ7nnB
5w3kOO7gsnbrsH4p0i75aBVyhshIUlCESLrwHuO/icSumIj+HQjgp8tepTsYNmCCwN2sHshf6sMR
5WXywAzgi/FcgKqKU83+zQsciaeVovj7KmgwdkmqnWBEMeFwt1OGl/BHqIuhuti1LzP3xA1VE19Q
/VC0iOdMgSIUACpnGV9Wa8Afz+clirVIrECKjdvejGhX/gByhaTI12YG/q0qCRryz+1iW7w7Qcph
GScyO4mlHbaORm4TbsekR7hO4gflUW4XuoH/MncokFm+h6OPdPXDiDM64iAtRlsCzr5gA2oxb9lv
hmjRR/EBTcix5XfodXT3GQEWGRmMxRdeP5lJ3I5paxdIMoWZKGdWPTofvj0UpCBo9+O+L/hUEk57
ND44HKPEGNTW2V0wS6R2To5cVZ5Lxu2YiVlW8B4MydMsa2xyClYpThHEV/WoeYQFifxD8Ii3ar9/
yhJ0SZHY/3FAAKZQWqtRB2YDx2H3HpGGtAz+lqX5A5DlAv/G9Xz1Dx2MB0Y50WiqJdrCX/qbCjdb
gwV4hA3JpB49gzDd9BY/vgQSxswzXIE8kzDAO3BeNDrP5iMZkpTxBtoN6UpER04DhnShlw9NcTf6
UYRavXqmxKd54h0O87Vo7ScOgyl8+hWkRv6zUuvhYpUuWfpG4wKCaoXSA/J+TgY+C1+GdS2kFKOx
acoZq14YOJ+oRYl1Nu38pBl2KBD96Vqse+L2KXMsmcx3j3lIG+G91sGKQRdtM2ExNOME16xBU07l
oL8fAPbGd/LrFw==
`protect end_protected
